# ------------------------------------------------------
#
#
#
#		RacyICs Memory Generator - RI MGene
#
#		DD/MM/YYYY Release Version
#		19/05/2016 Preliminary Release 1.0
#		25/08/2016 Software Release 1.0
#		09/09/2016 Software Release 1.0.1
#		28/09/2016 Software Release 1.0.2
#		05/10/2016 Software Release 1.0.3
#		06/10/2016 Software Release 1.0.4
#		01/12/2016 Software Release 1.0.5
#		01/12/2016 Software Release 1.0.6
#		09/02/2017 Software Release 1.0.7
#		17/02/2017 Software Release 1.0.8
#		09/03/2017 Software Release 1.0.9
#		10/08/2017 Software Release 1.0.10
#
#		Software Versions
#		RI MGene Memory Generator 1.0.10
#		RI MGene SRAM Explorer GUI 1.0
#		RI MGene Database Version 1.0.10082017
#
#		PDK Version
#		IHP SG13S rev1.0.2_a_150421
#		Generated on Tue Jun 14 11:44:36 2022		
#
# ------------------------------------------------------ 
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO RM_IHPSG13_1P_8192x32_c4_bm_bist
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN RM_IHPSG13_1P_8192x32_c4_bm_bist 0 0 ;
  SIZE 1520.16 BY 618.3 ;
  SYMMETRY X Y R90 ;
  PIN A_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 803.71 0 803.97 0.26 ;
    END
  END A_DIN[16]
  PIN A_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 716.19 0 716.45 0.26 ;
    END
  END A_DIN[15]
  PIN A_BIST_DIN[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 804.645 0 804.905 0.26 ;
    END
  END A_BIST_DIN[16]
  PIN A_BIST_DIN[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 715.255 0 715.515 0.26 ;
    END
  END A_BIST_DIN[15]
  PIN A_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 842.67 0 842.93 0.26 ;
    END
  END A_BM[16]
  PIN A_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 677.23 0 677.49 0.26 ;
    END
  END A_BM[15]
  PIN A_BIST_BM[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 841.14 0 841.4 0.26 ;
    END
  END A_BIST_BM[16]
  PIN A_BIST_BM[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 678.76 0 679.02 0.26 ;
    END
  END A_BIST_BM[15]
  PIN A_DOUT[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 825.485 0 825.745 0.26 ;
    END
  END A_DOUT[16]
  PIN A_DOUT[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 694.415 0 694.675 0.26 ;
    END
  END A_DOUT[15]
  PIN VSS!
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "vss VSS!" ;
    PORT
      LAYER Metal4 ;
        RECT 1496.23 0 1499.04 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1484.99 0 1487.8 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1473.75 0 1476.56 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1451.27 0 1454.08 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1440.03 0 1442.84 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1428.79 0 1431.6 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1406.31 0 1409.12 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1395.07 0 1397.88 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1383.83 0 1386.64 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1361.35 0 1364.16 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1350.11 0 1352.92 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1338.87 0 1341.68 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1316.39 0 1319.2 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1305.15 0 1307.96 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1293.91 0 1296.72 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1271.43 0 1274.24 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1260.19 0 1263 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1248.95 0 1251.76 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1226.47 0 1229.28 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1215.23 0 1218.04 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1203.99 0 1206.8 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1181.51 0 1184.32 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1170.27 0 1173.08 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1159.03 0 1161.84 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1136.55 0 1139.36 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1125.31 0 1128.12 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1114.07 0 1116.88 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1091.59 0 1094.4 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1080.35 0 1083.16 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1069.11 0 1071.92 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1046.63 0 1049.44 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1035.39 0 1038.2 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1024.15 0 1026.96 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1001.67 0 1004.48 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 990.43 0 993.24 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 979.19 0 982 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 956.71 0 959.52 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 945.47 0 948.28 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 934.23 0 937.04 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 911.75 0 914.56 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 900.51 0 903.32 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 889.27 0 892.08 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 866.79 0 869.6 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 855.55 0 858.36 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 844.31 0 847.12 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 821.83 0 824.64 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 810.59 0 813.4 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 799.35 0 802.16 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 776.7 0 779.51 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 766.4 0 769.21 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 750.95 0 753.76 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 740.65 0 743.46 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 718 0 720.81 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 706.76 0 709.57 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 695.52 0 698.33 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 673.04 0 675.85 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 661.8 0 664.61 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 650.56 0 653.37 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 628.08 0 630.89 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 616.84 0 619.65 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 605.6 0 608.41 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 583.12 0 585.93 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 571.88 0 574.69 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 560.64 0 563.45 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 538.16 0 540.97 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 526.92 0 529.73 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 515.68 0 518.49 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 493.2 0 496.01 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 481.96 0 484.77 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 470.72 0 473.53 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 448.24 0 451.05 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 437 0 439.81 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 425.76 0 428.57 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 403.28 0 406.09 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 392.04 0 394.85 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 380.8 0 383.61 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 358.32 0 361.13 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 347.08 0 349.89 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 335.84 0 338.65 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 313.36 0 316.17 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 302.12 0 304.93 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 290.88 0 293.69 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 268.4 0 271.21 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 257.16 0 259.97 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 245.92 0 248.73 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 223.44 0 226.25 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 212.2 0 215.01 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 200.96 0 203.77 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 178.48 0 181.29 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 167.24 0 170.05 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 156 0 158.81 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 133.52 0 136.33 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 122.28 0 125.09 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 111.04 0 113.85 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 88.56 0 91.37 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 77.32 0 80.13 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 66.08 0 68.89 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 43.6 0 46.41 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 32.36 0 35.17 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 21.12 0 23.93 618.3 ;
    END
  END VSS!
  PIN VDD!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vdd VDD!" ;
    PORT
      LAYER Metal4 ;
        RECT 1501.85 0 1504.66 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1490.61 0 1493.42 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1479.37 0 1482.18 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1456.89 0 1459.7 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1445.65 0 1448.46 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1434.41 0 1437.22 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1411.93 0 1414.74 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1400.69 0 1403.5 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1389.45 0 1392.26 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1366.97 0 1369.78 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1355.73 0 1358.54 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1344.49 0 1347.3 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1322.01 0 1324.82 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1310.77 0 1313.58 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1299.53 0 1302.34 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1277.05 0 1279.86 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1265.81 0 1268.62 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1254.57 0 1257.38 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1232.09 0 1234.9 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1220.85 0 1223.66 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1209.61 0 1212.42 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1187.13 0 1189.94 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1175.89 0 1178.7 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1164.65 0 1167.46 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1142.17 0 1144.98 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1130.93 0 1133.74 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1119.69 0 1122.5 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.21 0 1100.02 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1085.97 0 1088.78 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1074.73 0 1077.54 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1052.25 0 1055.06 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1041.01 0 1043.82 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1029.77 0 1032.58 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1007.29 0 1010.1 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 996.05 0 998.86 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 984.81 0 987.62 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 962.33 0 965.14 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 951.09 0 953.9 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 939.85 0 942.66 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 917.37 0 920.18 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 906.13 0 908.94 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 894.89 0 897.7 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 872.41 0 875.22 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 861.17 0 863.98 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 849.93 0 852.74 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 827.45 0 830.26 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 816.21 0 819.02 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 804.97 0 807.78 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 771.55 0 774.36 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 761.25 0 764.06 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 756.1 0 758.91 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 745.8 0 748.61 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 712.38 0 715.19 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 701.14 0 703.95 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 689.9 0 692.71 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 667.42 0 670.23 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 656.18 0 658.99 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 644.94 0 647.75 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 622.46 0 625.27 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 611.22 0 614.03 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 599.98 0 602.79 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 577.5 0 580.31 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 566.26 0 569.07 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.02 0 557.83 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 532.54 0 535.35 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 521.3 0 524.11 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 510.06 0 512.87 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 487.58 0 490.39 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 476.34 0 479.15 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 465.1 0 467.91 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 442.62 0 445.43 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 431.38 0 434.19 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 420.14 0 422.95 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 397.66 0 400.47 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 386.42 0 389.23 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.18 0 377.99 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.7 0 355.51 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 341.46 0 344.27 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.22 0 333.03 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 307.74 0 310.55 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 296.5 0 299.31 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.26 0 288.07 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.78 0 265.59 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 251.54 0 254.35 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.3 0 243.11 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 217.82 0 220.63 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206.58 0 209.39 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 195.34 0 198.15 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 0 175.67 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 0 164.43 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 0 153.19 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 0 130.71 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 0 119.47 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 0 108.23 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 0 85.75 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 0 74.51 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 0 63.27 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 0 40.79 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 0 29.55 30.425 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 0 18.31 30.425 ;
    END
  END VDD!
  PIN VDDARRAY!
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "vddarray VDDARRAY!" ;
    PORT
      LAYER Metal4 ;
        RECT 1501.85 37.065 1504.66 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1490.61 37.065 1493.42 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1479.37 37.065 1482.18 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1456.89 37.065 1459.7 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1445.65 37.065 1448.46 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1434.41 37.065 1437.22 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1411.93 37.065 1414.74 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1400.69 37.065 1403.5 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1389.45 37.065 1392.26 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1366.97 37.065 1369.78 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1355.73 37.065 1358.54 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1344.49 37.065 1347.3 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1322.01 37.065 1324.82 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1310.77 37.065 1313.58 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1299.53 37.065 1302.34 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1277.05 37.065 1279.86 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1265.81 37.065 1268.62 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1254.57 37.065 1257.38 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1232.09 37.065 1234.9 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1220.85 37.065 1223.66 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1209.61 37.065 1212.42 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1187.13 37.065 1189.94 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1175.89 37.065 1178.7 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1164.65 37.065 1167.46 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1142.17 37.065 1144.98 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1130.93 37.065 1133.74 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1119.69 37.065 1122.5 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.21 37.065 1100.02 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1085.97 37.065 1088.78 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1074.73 37.065 1077.54 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1052.25 37.065 1055.06 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1041.01 37.065 1043.82 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1029.77 37.065 1032.58 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1007.29 37.065 1010.1 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 996.05 37.065 998.86 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 984.81 37.065 987.62 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 962.33 37.065 965.14 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 951.09 37.065 953.9 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 939.85 37.065 942.66 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 917.37 37.065 920.18 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 906.13 37.065 908.94 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 894.89 37.065 897.7 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 872.41 37.065 875.22 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 861.17 37.065 863.98 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 849.93 37.065 852.74 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 827.45 37.065 830.26 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 816.21 37.065 819.02 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 804.97 37.065 807.78 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 712.38 37.065 715.19 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 701.14 37.065 703.95 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 689.9 37.065 692.71 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 667.42 37.065 670.23 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 656.18 37.065 658.99 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 644.94 37.065 647.75 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 622.46 37.065 625.27 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 611.22 37.065 614.03 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 599.98 37.065 602.79 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 577.5 37.065 580.31 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 566.26 37.065 569.07 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 555.02 37.065 557.83 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 532.54 37.065 535.35 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 521.3 37.065 524.11 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 510.06 37.065 512.87 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 487.58 37.065 490.39 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 476.34 37.065 479.15 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 465.1 37.065 467.91 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 442.62 37.065 445.43 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 431.38 37.065 434.19 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 420.14 37.065 422.95 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 397.66 37.065 400.47 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 386.42 37.065 389.23 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 375.18 37.065 377.99 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 352.7 37.065 355.51 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 341.46 37.065 344.27 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 330.22 37.065 333.03 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 307.74 37.065 310.55 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 296.5 37.065 299.31 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 285.26 37.065 288.07 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 262.78 37.065 265.59 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 251.54 37.065 254.35 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 240.3 37.065 243.11 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 217.82 37.065 220.63 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 206.58 37.065 209.39 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 195.34 37.065 198.15 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 172.86 37.065 175.67 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 161.62 37.065 164.43 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 150.38 37.065 153.19 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 127.9 37.065 130.71 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 116.66 37.065 119.47 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 105.42 37.065 108.23 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 82.94 37.065 85.75 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 71.7 37.065 74.51 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 60.46 37.065 63.27 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 37.98 37.065 40.79 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 26.74 37.065 29.55 618.3 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 15.5 37.065 18.31 618.3 ;
    END
  END VDDARRAY!
  PIN A_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 848.67 0 848.93 0.26 ;
    END
  END A_DIN[17]
  PIN A_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 671.23 0 671.49 0.26 ;
    END
  END A_DIN[14]
  PIN A_BIST_DIN[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 849.605 0 849.865 0.26 ;
    END
  END A_BIST_DIN[17]
  PIN A_BIST_DIN[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 670.295 0 670.555 0.26 ;
    END
  END A_BIST_DIN[14]
  PIN A_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 887.63 0 887.89 0.26 ;
    END
  END A_BM[17]
  PIN A_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 632.27 0 632.53 0.26 ;
    END
  END A_BM[14]
  PIN A_BIST_BM[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 886.1 0 886.36 0.26 ;
    END
  END A_BIST_BM[17]
  PIN A_BIST_BM[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 633.8 0 634.06 0.26 ;
    END
  END A_BIST_BM[14]
  PIN A_DOUT[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 870.445 0 870.705 0.26 ;
    END
  END A_DOUT[17]
  PIN A_DOUT[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 649.455 0 649.715 0.26 ;
    END
  END A_DOUT[14]
  PIN A_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 893.63 0 893.89 0.26 ;
    END
  END A_DIN[18]
  PIN A_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 626.27 0 626.53 0.26 ;
    END
  END A_DIN[13]
  PIN A_BIST_DIN[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 894.565 0 894.825 0.26 ;
    END
  END A_BIST_DIN[18]
  PIN A_BIST_DIN[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 625.335 0 625.595 0.26 ;
    END
  END A_BIST_DIN[13]
  PIN A_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 932.59 0 932.85 0.26 ;
    END
  END A_BM[18]
  PIN A_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 587.31 0 587.57 0.26 ;
    END
  END A_BM[13]
  PIN A_BIST_BM[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 931.06 0 931.32 0.26 ;
    END
  END A_BIST_BM[18]
  PIN A_BIST_BM[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 588.84 0 589.1 0.26 ;
    END
  END A_BIST_BM[13]
  PIN A_DOUT[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 915.405 0 915.665 0.26 ;
    END
  END A_DOUT[18]
  PIN A_DOUT[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 604.495 0 604.755 0.26 ;
    END
  END A_DOUT[13]
  PIN A_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 938.59 0 938.85 0.26 ;
    END
  END A_DIN[19]
  PIN A_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 581.31 0 581.57 0.26 ;
    END
  END A_DIN[12]
  PIN A_BIST_DIN[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 939.525 0 939.785 0.26 ;
    END
  END A_BIST_DIN[19]
  PIN A_BIST_DIN[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 580.375 0 580.635 0.26 ;
    END
  END A_BIST_DIN[12]
  PIN A_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 977.55 0 977.81 0.26 ;
    END
  END A_BM[19]
  PIN A_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 542.35 0 542.61 0.26 ;
    END
  END A_BM[12]
  PIN A_BIST_BM[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 976.02 0 976.28 0.26 ;
    END
  END A_BIST_BM[19]
  PIN A_BIST_BM[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 543.88 0 544.14 0.26 ;
    END
  END A_BIST_BM[12]
  PIN A_DOUT[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 960.365 0 960.625 0.26 ;
    END
  END A_DOUT[19]
  PIN A_DOUT[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 559.535 0 559.795 0.26 ;
    END
  END A_DOUT[12]
  PIN A_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 983.55 0 983.81 0.26 ;
    END
  END A_DIN[20]
  PIN A_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 536.35 0 536.61 0.26 ;
    END
  END A_DIN[11]
  PIN A_BIST_DIN[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 984.485 0 984.745 0.26 ;
    END
  END A_BIST_DIN[20]
  PIN A_BIST_DIN[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 535.415 0 535.675 0.26 ;
    END
  END A_BIST_DIN[11]
  PIN A_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1022.51 0 1022.77 0.26 ;
    END
  END A_BM[20]
  PIN A_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 497.39 0 497.65 0.26 ;
    END
  END A_BM[11]
  PIN A_BIST_BM[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1020.98 0 1021.24 0.26 ;
    END
  END A_BIST_BM[20]
  PIN A_BIST_BM[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 498.92 0 499.18 0.26 ;
    END
  END A_BIST_BM[11]
  PIN A_DOUT[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1005.325 0 1005.585 0.26 ;
    END
  END A_DOUT[20]
  PIN A_DOUT[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 514.575 0 514.835 0.26 ;
    END
  END A_DOUT[11]
  PIN A_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1028.51 0 1028.77 0.26 ;
    END
  END A_DIN[21]
  PIN A_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 491.39 0 491.65 0.26 ;
    END
  END A_DIN[10]
  PIN A_BIST_DIN[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1029.445 0 1029.705 0.26 ;
    END
  END A_BIST_DIN[21]
  PIN A_BIST_DIN[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 490.455 0 490.715 0.26 ;
    END
  END A_BIST_DIN[10]
  PIN A_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1067.47 0 1067.73 0.26 ;
    END
  END A_BM[21]
  PIN A_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 452.43 0 452.69 0.26 ;
    END
  END A_BM[10]
  PIN A_BIST_BM[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1065.94 0 1066.2 0.26 ;
    END
  END A_BIST_BM[21]
  PIN A_BIST_BM[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 453.96 0 454.22 0.26 ;
    END
  END A_BIST_BM[10]
  PIN A_DOUT[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1050.285 0 1050.545 0.26 ;
    END
  END A_DOUT[21]
  PIN A_DOUT[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 469.615 0 469.875 0.26 ;
    END
  END A_DOUT[10]
  PIN A_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1073.47 0 1073.73 0.26 ;
    END
  END A_DIN[22]
  PIN A_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 446.43 0 446.69 0.26 ;
    END
  END A_DIN[9]
  PIN A_BIST_DIN[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1074.405 0 1074.665 0.26 ;
    END
  END A_BIST_DIN[22]
  PIN A_BIST_DIN[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 445.495 0 445.755 0.26 ;
    END
  END A_BIST_DIN[9]
  PIN A_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1112.43 0 1112.69 0.26 ;
    END
  END A_BM[22]
  PIN A_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 407.47 0 407.73 0.26 ;
    END
  END A_BM[9]
  PIN A_BIST_BM[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1110.9 0 1111.16 0.26 ;
    END
  END A_BIST_BM[22]
  PIN A_BIST_BM[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 409 0 409.26 0.26 ;
    END
  END A_BIST_BM[9]
  PIN A_DOUT[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1095.245 0 1095.505 0.26 ;
    END
  END A_DOUT[22]
  PIN A_DOUT[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 424.655 0 424.915 0.26 ;
    END
  END A_DOUT[9]
  PIN A_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1118.43 0 1118.69 0.26 ;
    END
  END A_DIN[23]
  PIN A_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 401.47 0 401.73 0.26 ;
    END
  END A_DIN[8]
  PIN A_BIST_DIN[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1119.365 0 1119.625 0.26 ;
    END
  END A_BIST_DIN[23]
  PIN A_BIST_DIN[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 400.535 0 400.795 0.26 ;
    END
  END A_BIST_DIN[8]
  PIN A_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1157.39 0 1157.65 0.26 ;
    END
  END A_BM[23]
  PIN A_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 362.51 0 362.77 0.26 ;
    END
  END A_BM[8]
  PIN A_BIST_BM[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1155.86 0 1156.12 0.26 ;
    END
  END A_BIST_BM[23]
  PIN A_BIST_BM[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 364.04 0 364.3 0.26 ;
    END
  END A_BIST_BM[8]
  PIN A_DOUT[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1140.205 0 1140.465 0.26 ;
    END
  END A_DOUT[23]
  PIN A_DOUT[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 379.695 0 379.955 0.26 ;
    END
  END A_DOUT[8]
  PIN A_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1163.39 0 1163.65 0.26 ;
    END
  END A_DIN[24]
  PIN A_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 356.51 0 356.77 0.26 ;
    END
  END A_DIN[7]
  PIN A_BIST_DIN[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1164.325 0 1164.585 0.26 ;
    END
  END A_BIST_DIN[24]
  PIN A_BIST_DIN[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 355.575 0 355.835 0.26 ;
    END
  END A_BIST_DIN[7]
  PIN A_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1202.35 0 1202.61 0.26 ;
    END
  END A_BM[24]
  PIN A_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 317.55 0 317.81 0.26 ;
    END
  END A_BM[7]
  PIN A_BIST_BM[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1200.82 0 1201.08 0.26 ;
    END
  END A_BIST_BM[24]
  PIN A_BIST_BM[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 319.08 0 319.34 0.26 ;
    END
  END A_BIST_BM[7]
  PIN A_DOUT[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1185.165 0 1185.425 0.26 ;
    END
  END A_DOUT[24]
  PIN A_DOUT[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 334.735 0 334.995 0.26 ;
    END
  END A_DOUT[7]
  PIN A_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1208.35 0 1208.61 0.26 ;
    END
  END A_DIN[25]
  PIN A_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 311.55 0 311.81 0.26 ;
    END
  END A_DIN[6]
  PIN A_BIST_DIN[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1209.285 0 1209.545 0.26 ;
    END
  END A_BIST_DIN[25]
  PIN A_BIST_DIN[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 310.615 0 310.875 0.26 ;
    END
  END A_BIST_DIN[6]
  PIN A_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1247.31 0 1247.57 0.26 ;
    END
  END A_BM[25]
  PIN A_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 272.59 0 272.85 0.26 ;
    END
  END A_BM[6]
  PIN A_BIST_BM[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1245.78 0 1246.04 0.26 ;
    END
  END A_BIST_BM[25]
  PIN A_BIST_BM[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 274.12 0 274.38 0.26 ;
    END
  END A_BIST_BM[6]
  PIN A_DOUT[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1230.125 0 1230.385 0.26 ;
    END
  END A_DOUT[25]
  PIN A_DOUT[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 289.775 0 290.035 0.26 ;
    END
  END A_DOUT[6]
  PIN A_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1253.31 0 1253.57 0.26 ;
    END
  END A_DIN[26]
  PIN A_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 266.59 0 266.85 0.26 ;
    END
  END A_DIN[5]
  PIN A_BIST_DIN[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1254.245 0 1254.505 0.26 ;
    END
  END A_BIST_DIN[26]
  PIN A_BIST_DIN[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 265.655 0 265.915 0.26 ;
    END
  END A_BIST_DIN[5]
  PIN A_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1292.27 0 1292.53 0.26 ;
    END
  END A_BM[26]
  PIN A_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 227.63 0 227.89 0.26 ;
    END
  END A_BM[5]
  PIN A_BIST_BM[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1290.74 0 1291 0.26 ;
    END
  END A_BIST_BM[26]
  PIN A_BIST_BM[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 229.16 0 229.42 0.26 ;
    END
  END A_BIST_BM[5]
  PIN A_DOUT[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1275.085 0 1275.345 0.26 ;
    END
  END A_DOUT[26]
  PIN A_DOUT[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 244.815 0 245.075 0.26 ;
    END
  END A_DOUT[5]
  PIN A_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1298.27 0 1298.53 0.26 ;
    END
  END A_DIN[27]
  PIN A_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 221.63 0 221.89 0.26 ;
    END
  END A_DIN[4]
  PIN A_BIST_DIN[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1299.205 0 1299.465 0.26 ;
    END
  END A_BIST_DIN[27]
  PIN A_BIST_DIN[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 220.695 0 220.955 0.26 ;
    END
  END A_BIST_DIN[4]
  PIN A_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1337.23 0 1337.49 0.26 ;
    END
  END A_BM[27]
  PIN A_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 182.67 0 182.93 0.26 ;
    END
  END A_BM[4]
  PIN A_BIST_BM[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1335.7 0 1335.96 0.26 ;
    END
  END A_BIST_BM[27]
  PIN A_BIST_BM[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 184.2 0 184.46 0.26 ;
    END
  END A_BIST_BM[4]
  PIN A_DOUT[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1320.045 0 1320.305 0.26 ;
    END
  END A_DOUT[27]
  PIN A_DOUT[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 199.855 0 200.115 0.26 ;
    END
  END A_DOUT[4]
  PIN A_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1343.23 0 1343.49 0.26 ;
    END
  END A_DIN[28]
  PIN A_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 176.67 0 176.93 0.26 ;
    END
  END A_DIN[3]
  PIN A_BIST_DIN[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1344.165 0 1344.425 0.26 ;
    END
  END A_BIST_DIN[28]
  PIN A_BIST_DIN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 175.735 0 175.995 0.26 ;
    END
  END A_BIST_DIN[3]
  PIN A_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1382.19 0 1382.45 0.26 ;
    END
  END A_BM[28]
  PIN A_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 137.71 0 137.97 0.26 ;
    END
  END A_BM[3]
  PIN A_BIST_BM[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1380.66 0 1380.92 0.26 ;
    END
  END A_BIST_BM[28]
  PIN A_BIST_BM[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 139.24 0 139.5 0.26 ;
    END
  END A_BIST_BM[3]
  PIN A_DOUT[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1365.005 0 1365.265 0.26 ;
    END
  END A_DOUT[28]
  PIN A_DOUT[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 154.895 0 155.155 0.26 ;
    END
  END A_DOUT[3]
  PIN A_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1388.19 0 1388.45 0.26 ;
    END
  END A_DIN[29]
  PIN A_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 131.71 0 131.97 0.26 ;
    END
  END A_DIN[2]
  PIN A_BIST_DIN[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1389.125 0 1389.385 0.26 ;
    END
  END A_BIST_DIN[29]
  PIN A_BIST_DIN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 130.775 0 131.035 0.26 ;
    END
  END A_BIST_DIN[2]
  PIN A_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1427.15 0 1427.41 0.26 ;
    END
  END A_BM[29]
  PIN A_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 92.75 0 93.01 0.26 ;
    END
  END A_BM[2]
  PIN A_BIST_BM[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1425.62 0 1425.88 0.26 ;
    END
  END A_BIST_BM[29]
  PIN A_BIST_BM[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 94.28 0 94.54 0.26 ;
    END
  END A_BIST_BM[2]
  PIN A_DOUT[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1409.965 0 1410.225 0.26 ;
    END
  END A_DOUT[29]
  PIN A_DOUT[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 109.935 0 110.195 0.26 ;
    END
  END A_DOUT[2]
  PIN A_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1433.15 0 1433.41 0.26 ;
    END
  END A_DIN[30]
  PIN A_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 86.75 0 87.01 0.26 ;
    END
  END A_DIN[1]
  PIN A_BIST_DIN[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1434.085 0 1434.345 0.26 ;
    END
  END A_BIST_DIN[30]
  PIN A_BIST_DIN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 85.815 0 86.075 0.26 ;
    END
  END A_BIST_DIN[1]
  PIN A_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1472.11 0 1472.37 0.26 ;
    END
  END A_BM[30]
  PIN A_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 47.79 0 48.05 0.26 ;
    END
  END A_BM[1]
  PIN A_BIST_BM[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1470.58 0 1470.84 0.26 ;
    END
  END A_BIST_BM[30]
  PIN A_BIST_BM[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 49.32 0 49.58 0.26 ;
    END
  END A_BIST_BM[1]
  PIN A_DOUT[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1454.925 0 1455.185 0.26 ;
    END
  END A_DOUT[30]
  PIN A_DOUT[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 64.975 0 65.235 0.26 ;
    END
  END A_DOUT[1]
  PIN A_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1478.11 0 1478.37 0.26 ;
    END
  END A_DIN[31]
  PIN A_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 41.79 0 42.05 0.26 ;
    END
  END A_DIN[0]
  PIN A_BIST_DIN[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1479.045 0 1479.305 0.26 ;
    END
  END A_BIST_DIN[31]
  PIN A_BIST_DIN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0394 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 16.038835 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 40.855 0 41.115 0.26 ;
    END
  END A_BIST_DIN[0]
  PIN A_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1517.07 0 1517.33 0.26 ;
    END
  END A_BM[31]
  PIN A_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 2.83 0 3.09 0.26 ;
    END
  END A_BM[0]
  PIN A_BIST_BM[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1515.54 0 1515.8 0.26 ;
    END
  END A_BIST_BM[31]
  PIN A_BIST_BM[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8847 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 15.268608 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 4.36 0 4.62 0.26 ;
    END
  END A_BIST_BM[0]
  PIN A_DOUT[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 1499.885 0 1500.145 0.26 ;
    END
  END A_DOUT[31]
  PIN A_DOUT[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5834 LAYER Metal2 ;
    ANTENNADIFFAREA 0.988 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 20.015 0 20.275 0.26 ;
    END
  END A_DOUT[0]
  PIN A_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.7171 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 34.349515 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 756.28 0 756.54 0.26 ;
    END
  END A_ADDR[0]
  PIN A_BIST_ADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5127 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 38.31068 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 760.87 0 761.13 0.26 ;
    END
  END A_BIST_ADDR[0]
  PIN A_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.59 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 28.783172 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 755.77 0 756.03 0.26 ;
    END
  END A_ADDR[1]
  PIN A_BIST_ADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3856 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 32.744337 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 760.36 0 760.62 0.26 ;
    END
  END A_BIST_ADDR[1]
  PIN A_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4519 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 33.029126 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 741.49 0 741.75 0.26 ;
    END
  END A_ADDR[2]
  PIN A_BIST_ADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1867 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 31.708738 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 743.02 0 743.28 0.26 ;
    END
  END A_BIST_ADDR[2]
  PIN A_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0947 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.2684 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 8.671148 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 746.08 0 746.34 0.26 ;
    END
  END A_ADDR[3]
  PIN A_BIST_ADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4395 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0542 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 10.866816 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 746.59 0 746.85 0.26 ;
    END
  END A_BIST_ADDR[3]
  PIN A_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5246 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.415982 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 763.93 0 764.19 0.26 ;
    END
  END A_ADDR[4]
  PIN A_BIST_ADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.0962 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 7.813791 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 764.44 0 764.7 0.26 ;
    END
  END A_BIST_ADDR[4]
  PIN A_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.8367 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 20.927558 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 762.91 0 763.17 0.26 ;
    END
  END A_ADDR[5]
  PIN A_BIST_ADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4487 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 3.5175 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 19.869057 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 763.42 0 763.68 0.26 ;
    END
  END A_BIST_ADDR[5]
  PIN A_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.0139 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 50.763754 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 766.48 0 766.74 0.26 ;
    END
  END A_ADDR[6]
  PIN A_BIST_ADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.7487 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 49.443366 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 765.97 0 766.23 0.26 ;
    END
  END A_BIST_ADDR[6]
  PIN A_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.7429 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 59.372168 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 765.46 0 765.72 0.26 ;
    END
  END A_ADDR[7]
  PIN A_BIST_ADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.4777 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 58.05178 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 764.95 0 765.21 0.26 ;
    END
  END A_BIST_ADDR[7]
  PIN A_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.7685 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 44.563107 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 744.04 0 744.3 0.26 ;
    END
  END A_ADDR[8]
  PIN A_BIST_ADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.4931 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.191934 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 744.55 0 744.81 0.26 ;
    END
  END A_BIST_ADDR[8]
  PIN A_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.2323 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 51.851133 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 745.06 0 745.32 0.26 ;
    END
  END A_ADDR[9]
  PIN A_BIST_ADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.9671 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 50.530744 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 745.57 0 745.83 0.26 ;
    END
  END A_BIST_ADDR[9]
  PIN A_ADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9183 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.5897 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.740105 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 774.13 0 774.39 0.26 ;
    END
  END A_ADDR[10]
  PIN A_BIST_ADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.9183 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 1.3755 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal3 ;
      ANTENNAMAXAREACAR 9.204381 LAYER Metal3 ;
    PORT
      LAYER Metal2 ;
        RECT 774.64 0 774.9 0.26 ;
    END
  END A_BIST_ADDR[10]
  PIN A_ADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.6097 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 53.730147 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 769.03 0 769.29 0.26 ;
    END
  END A_ADDR[11]
  PIN A_BIST_ADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.3547 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 52.460543 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 769.54 0 769.8 0.26 ;
    END
  END A_BIST_ADDR[11]
  PIN A_ADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6359 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.902913 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 766.99 0 767.25 0.26 ;
    END
  END A_ADDR[12]
  PIN A_BIST_ADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.6359 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 43.902913 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 767.5 0 767.76 0.26 ;
    END
  END A_BIST_ADDR[12]
  PIN A_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8707 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 10.220065 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 754.24 0 754.5 0.26 ;
    END
  END A_CLK
  PIN A_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.81105 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 9.923077 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 757.81 0 758.07 0.26 ;
    END
  END A_REN
  PIN A_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7007 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.394822 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 757.3 0 757.56 0.26 ;
    END
  END A_WEN
  PIN A_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8407 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 5.09186 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 754.75 0 755.01 0.26 ;
    END
  END A_MEN
  PIN A_DLY
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.874 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3367 LAYER Metal2 ;
      ANTENNAMAXAREACAR 12.046332 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 776.17 0 776.43 0.26 ;
    END
  END A_DLY
  PIN A_BIST_EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8031 LAYER Metal2 ;
    ANTENNAPARTIALMETALAREA 405.14255 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER Via2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.43 LAYER Metal2 ;
      ANTENNAGATEAREA 28.9575 LAYER Metal3 ;
      ANTENNAMAXAREACAR 1.686364 LAYER Metal2 ;
      ANTENNAMAXAREACAR 19.644028 LAYER Metal3 ;
      ANTENNAMAXCUTCAR 0.151469 LAYER Via2 ;
    PORT
      LAYER Metal2 ;
        RECT 756.79 0 757.05 0.26 ;
    END
  END A_BIST_EN
  PIN A_BIST_CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9799 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 11.079661 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 752.71 0 752.97 0.26 ;
    END
  END A_BIST_CLK
  PIN A_BIST_REN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9279 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 10.820762 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 759.34 0 759.6 0.26 ;
    END
  END A_BIST_REN
  PIN A_BIST_WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7211 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.812298 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 758.83 0 759.09 0.26 ;
    END
  END A_BIST_WEN
  PIN A_BIST_MEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7137 LAYER Metal2 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20085 LAYER Metal2 ;
      ANTENNAMAXAREACAR 4.775454 LAYER Metal2 ;
    PORT
      LAYER Metal2 ;
        RECT 753.22 0 753.48 0.26 ;
    END
  END A_BIST_MEN
  OBS
    LAYER Metal1 ;
      RECT 0 0 1520.16 618.3 ;
    LAYER Metal2 ;
      RECT 0.105 37.065 0.305 618.275 ;
      RECT 1.1 617.545 1.3 618.275 ;
      RECT 1.92 617.545 2.12 618.275 ;
      RECT 2.415 617.545 2.615 618.275 ;
      RECT 2.83 0.52 3.09 7.94 ;
      RECT 2.915 617.545 3.115 618.275 ;
      RECT 3.415 617.545 3.615 618.275 ;
      RECT 3.91 617.545 4.11 618.275 ;
      RECT 4.36 0.52 4.62 10.655 ;
      RECT 5.225 0.17 5.995 0.43 ;
      RECT 5.735 0.17 5.995 11.38 ;
      RECT 5.225 0.17 5.485 16.7 ;
      RECT 4.73 617.545 4.93 618.275 ;
      RECT 5.225 617.545 5.425 618.275 ;
      RECT 5.725 617.545 5.925 618.275 ;
      RECT 6.225 617.545 6.425 618.275 ;
      RECT 6.72 617.545 6.92 618.275 ;
      RECT 7.54 617.545 7.74 618.275 ;
      RECT 8.795 0.17 9.565 0.43 ;
      RECT 9.305 0.17 9.565 8.7 ;
      RECT 8.795 0.17 9.055 16.7 ;
      RECT 8.035 617.545 8.235 618.275 ;
      RECT 8.535 617.545 8.735 618.275 ;
      RECT 9.035 617.545 9.235 618.275 ;
      RECT 9.53 617.545 9.73 618.275 ;
      RECT 9.815 0.3 10.075 4.63 ;
      RECT 10.35 617.545 10.55 618.275 ;
      RECT 10.835 0.17 11.605 0.43 ;
      RECT 11.345 0.17 11.605 8.7 ;
      RECT 10.835 0.17 11.095 16.7 ;
      RECT 10.325 0.3 10.585 4.63 ;
      RECT 10.845 617.545 11.045 618.275 ;
      RECT 11.345 617.545 11.545 618.275 ;
      RECT 11.845 617.545 12.045 618.275 ;
      RECT 12.34 617.545 12.54 618.275 ;
      RECT 13.16 617.545 13.36 618.275 ;
      RECT 13.655 617.545 13.855 618.275 ;
      RECT 14.155 617.545 14.355 618.275 ;
      RECT 14.655 617.545 14.855 618.275 ;
      RECT 15.15 617.545 15.35 618.275 ;
      RECT 15.97 617.545 16.17 618.275 ;
      RECT 16.465 617.545 16.665 618.275 ;
      RECT 16.965 617.545 17.165 618.275 ;
      RECT 17.465 617.545 17.665 618.275 ;
      RECT 17.565 0.3 17.825 4.63 ;
      RECT 18.585 0.165 19.355 0.425 ;
      RECT 18.585 0.165 18.845 8.825 ;
      RECT 19.095 0.165 19.355 8.825 ;
      RECT 17.96 617.545 18.16 618.275 ;
      RECT 18.075 0.3 18.335 4.63 ;
      RECT 18.78 617.545 18.98 618.275 ;
      RECT 19.275 617.545 19.475 618.275 ;
      RECT 19.775 617.545 19.975 618.275 ;
      RECT 20.015 0.52 20.275 4.5 ;
      RECT 20.275 617.545 20.475 618.275 ;
      RECT 20.77 617.545 20.97 618.275 ;
      RECT 21.59 617.545 21.79 618.275 ;
      RECT 22.085 617.545 22.285 618.275 ;
      RECT 22.585 617.545 22.785 618.275 ;
      RECT 23.085 617.545 23.285 618.275 ;
      RECT 23.58 617.545 23.78 618.275 ;
      RECT 24.4 617.545 24.6 618.275 ;
      RECT 24.895 617.545 25.095 618.275 ;
      RECT 25.395 617.545 25.595 618.275 ;
      RECT 25.895 617.545 26.095 618.275 ;
      RECT 26.39 617.545 26.59 618.275 ;
      RECT 27.21 617.545 27.41 618.275 ;
      RECT 27.705 617.545 27.905 618.275 ;
      RECT 28.205 617.545 28.405 618.275 ;
      RECT 28.705 617.545 28.905 618.275 ;
      RECT 29.2 617.545 29.4 618.275 ;
      RECT 30.02 617.545 30.22 618.275 ;
      RECT 30.515 617.545 30.715 618.275 ;
      RECT 31.015 617.545 31.215 618.275 ;
      RECT 31.515 617.545 31.715 618.275 ;
      RECT 32.01 617.545 32.21 618.275 ;
      RECT 32.83 617.545 33.03 618.275 ;
      RECT 33.785 0.16 34.555 0.42 ;
      RECT 34.295 0.16 34.555 4.63 ;
      RECT 33.785 0.16 34.045 8.82 ;
      RECT 33.325 617.545 33.525 618.275 ;
      RECT 33.825 617.545 34.025 618.275 ;
      RECT 34.325 617.545 34.525 618.275 ;
      RECT 34.82 617.545 35.02 618.275 ;
      RECT 34.805 0.3 35.065 4.63 ;
      RECT 35.315 0.3 35.575 4.63 ;
      RECT 35.64 617.545 35.84 618.275 ;
      RECT 36.135 617.545 36.335 618.275 ;
      RECT 36.635 617.545 36.835 618.275 ;
      RECT 38.32 0.16 39.09 0.42 ;
      RECT 38.32 0.16 38.58 8.82 ;
      RECT 38.83 0.16 39.09 8.82 ;
      RECT 37.135 617.545 37.335 618.275 ;
      RECT 37.63 617.545 37.83 618.275 ;
      RECT 38.45 617.545 38.65 618.275 ;
      RECT 38.945 617.545 39.145 618.275 ;
      RECT 39.34 0.3 39.6 4.63 ;
      RECT 39.445 617.545 39.645 618.275 ;
      RECT 39.85 0.3 40.11 4.63 ;
      RECT 39.945 617.545 40.145 618.275 ;
      RECT 40.44 617.545 40.64 618.275 ;
      RECT 40.855 0.52 41.115 10.655 ;
      RECT 41.26 617.545 41.46 618.275 ;
      RECT 41.755 617.545 41.955 618.275 ;
      RECT 41.79 0.52 42.05 4.5 ;
      RECT 42.255 617.545 42.455 618.275 ;
      RECT 42.755 617.545 42.955 618.275 ;
      RECT 43.25 617.545 43.45 618.275 ;
      RECT 44.495 0.165 45.265 0.425 ;
      RECT 44.495 0.165 44.755 8.825 ;
      RECT 45.005 0.165 45.265 8.825 ;
      RECT 44.07 617.545 44.27 618.275 ;
      RECT 44.565 617.545 44.765 618.275 ;
      RECT 45.065 617.545 45.265 618.275 ;
      RECT 45.565 617.545 45.765 618.275 ;
      RECT 45.515 0.3 45.775 4.63 ;
      RECT 46.06 617.545 46.26 618.275 ;
      RECT 46.025 0.3 46.285 8.23 ;
      RECT 46.88 617.545 47.08 618.275 ;
      RECT 47.375 617.545 47.575 618.275 ;
      RECT 47.79 0.52 48.05 7.94 ;
      RECT 47.875 617.545 48.075 618.275 ;
      RECT 48.375 617.545 48.575 618.275 ;
      RECT 48.87 617.545 49.07 618.275 ;
      RECT 49.32 0.52 49.58 10.655 ;
      RECT 50.185 0.17 50.955 0.43 ;
      RECT 50.695 0.17 50.955 11.38 ;
      RECT 50.185 0.17 50.445 16.7 ;
      RECT 49.69 617.545 49.89 618.275 ;
      RECT 50.185 617.545 50.385 618.275 ;
      RECT 50.685 617.545 50.885 618.275 ;
      RECT 51.185 617.545 51.385 618.275 ;
      RECT 51.68 617.545 51.88 618.275 ;
      RECT 52.5 617.545 52.7 618.275 ;
      RECT 53.755 0.17 54.525 0.43 ;
      RECT 54.265 0.17 54.525 8.7 ;
      RECT 53.755 0.17 54.015 16.7 ;
      RECT 52.995 617.545 53.195 618.275 ;
      RECT 53.495 617.545 53.695 618.275 ;
      RECT 53.995 617.545 54.195 618.275 ;
      RECT 54.49 617.545 54.69 618.275 ;
      RECT 54.775 0.3 55.035 4.63 ;
      RECT 55.31 617.545 55.51 618.275 ;
      RECT 55.795 0.17 56.565 0.43 ;
      RECT 56.305 0.17 56.565 8.7 ;
      RECT 55.795 0.17 56.055 16.7 ;
      RECT 55.285 0.3 55.545 4.63 ;
      RECT 55.805 617.545 56.005 618.275 ;
      RECT 56.305 617.545 56.505 618.275 ;
      RECT 56.805 617.545 57.005 618.275 ;
      RECT 57.3 617.545 57.5 618.275 ;
      RECT 58.12 617.545 58.32 618.275 ;
      RECT 58.615 617.545 58.815 618.275 ;
      RECT 59.115 617.545 59.315 618.275 ;
      RECT 59.615 617.545 59.815 618.275 ;
      RECT 60.11 617.545 60.31 618.275 ;
      RECT 60.93 617.545 61.13 618.275 ;
      RECT 61.425 617.545 61.625 618.275 ;
      RECT 61.925 617.545 62.125 618.275 ;
      RECT 62.425 617.545 62.625 618.275 ;
      RECT 62.525 0.3 62.785 4.63 ;
      RECT 63.545 0.165 64.315 0.425 ;
      RECT 63.545 0.165 63.805 8.825 ;
      RECT 64.055 0.165 64.315 8.825 ;
      RECT 62.92 617.545 63.12 618.275 ;
      RECT 63.035 0.3 63.295 4.63 ;
      RECT 63.74 617.545 63.94 618.275 ;
      RECT 64.235 617.545 64.435 618.275 ;
      RECT 64.735 617.545 64.935 618.275 ;
      RECT 64.975 0.52 65.235 4.5 ;
      RECT 65.235 617.545 65.435 618.275 ;
      RECT 65.73 617.545 65.93 618.275 ;
      RECT 66.55 617.545 66.75 618.275 ;
      RECT 67.045 617.545 67.245 618.275 ;
      RECT 67.545 617.545 67.745 618.275 ;
      RECT 68.045 617.545 68.245 618.275 ;
      RECT 68.54 617.545 68.74 618.275 ;
      RECT 69.36 617.545 69.56 618.275 ;
      RECT 69.855 617.545 70.055 618.275 ;
      RECT 70.355 617.545 70.555 618.275 ;
      RECT 70.855 617.545 71.055 618.275 ;
      RECT 71.35 617.545 71.55 618.275 ;
      RECT 72.17 617.545 72.37 618.275 ;
      RECT 72.665 617.545 72.865 618.275 ;
      RECT 73.165 617.545 73.365 618.275 ;
      RECT 73.665 617.545 73.865 618.275 ;
      RECT 74.16 617.545 74.36 618.275 ;
      RECT 74.98 617.545 75.18 618.275 ;
      RECT 75.475 617.545 75.675 618.275 ;
      RECT 75.975 617.545 76.175 618.275 ;
      RECT 76.475 617.545 76.675 618.275 ;
      RECT 76.97 617.545 77.17 618.275 ;
      RECT 77.79 617.545 77.99 618.275 ;
      RECT 78.745 0.16 79.515 0.42 ;
      RECT 79.255 0.16 79.515 4.63 ;
      RECT 78.745 0.16 79.005 8.82 ;
      RECT 78.285 617.545 78.485 618.275 ;
      RECT 78.785 617.545 78.985 618.275 ;
      RECT 79.285 617.545 79.485 618.275 ;
      RECT 79.78 617.545 79.98 618.275 ;
      RECT 79.765 0.3 80.025 4.63 ;
      RECT 80.275 0.3 80.535 4.63 ;
      RECT 80.6 617.545 80.8 618.275 ;
      RECT 81.095 617.545 81.295 618.275 ;
      RECT 81.595 617.545 81.795 618.275 ;
      RECT 83.28 0.16 84.05 0.42 ;
      RECT 83.28 0.16 83.54 8.82 ;
      RECT 83.79 0.16 84.05 8.82 ;
      RECT 82.095 617.545 82.295 618.275 ;
      RECT 82.59 617.545 82.79 618.275 ;
      RECT 83.41 617.545 83.61 618.275 ;
      RECT 83.905 617.545 84.105 618.275 ;
      RECT 84.3 0.3 84.56 4.63 ;
      RECT 84.405 617.545 84.605 618.275 ;
      RECT 84.81 0.3 85.07 4.63 ;
      RECT 84.905 617.545 85.105 618.275 ;
      RECT 85.4 617.545 85.6 618.275 ;
      RECT 85.815 0.52 86.075 10.655 ;
      RECT 86.22 617.545 86.42 618.275 ;
      RECT 86.715 617.545 86.915 618.275 ;
      RECT 86.75 0.52 87.01 4.5 ;
      RECT 87.215 617.545 87.415 618.275 ;
      RECT 87.715 617.545 87.915 618.275 ;
      RECT 88.21 617.545 88.41 618.275 ;
      RECT 89.455 0.165 90.225 0.425 ;
      RECT 89.455 0.165 89.715 8.825 ;
      RECT 89.965 0.165 90.225 8.825 ;
      RECT 89.03 617.545 89.23 618.275 ;
      RECT 89.525 617.545 89.725 618.275 ;
      RECT 90.025 617.545 90.225 618.275 ;
      RECT 90.525 617.545 90.725 618.275 ;
      RECT 90.475 0.3 90.735 4.63 ;
      RECT 91.02 617.545 91.22 618.275 ;
      RECT 90.985 0.3 91.245 8.23 ;
      RECT 91.84 617.545 92.04 618.275 ;
      RECT 92.335 617.545 92.535 618.275 ;
      RECT 92.75 0.52 93.01 7.94 ;
      RECT 92.835 617.545 93.035 618.275 ;
      RECT 93.335 617.545 93.535 618.275 ;
      RECT 93.83 617.545 94.03 618.275 ;
      RECT 94.28 0.52 94.54 10.655 ;
      RECT 95.145 0.17 95.915 0.43 ;
      RECT 95.655 0.17 95.915 11.38 ;
      RECT 95.145 0.17 95.405 16.7 ;
      RECT 94.65 617.545 94.85 618.275 ;
      RECT 95.145 617.545 95.345 618.275 ;
      RECT 95.645 617.545 95.845 618.275 ;
      RECT 96.145 617.545 96.345 618.275 ;
      RECT 96.64 617.545 96.84 618.275 ;
      RECT 97.46 617.545 97.66 618.275 ;
      RECT 98.715 0.17 99.485 0.43 ;
      RECT 99.225 0.17 99.485 8.7 ;
      RECT 98.715 0.17 98.975 16.7 ;
      RECT 97.955 617.545 98.155 618.275 ;
      RECT 98.455 617.545 98.655 618.275 ;
      RECT 98.955 617.545 99.155 618.275 ;
      RECT 99.45 617.545 99.65 618.275 ;
      RECT 99.735 0.3 99.995 4.63 ;
      RECT 100.27 617.545 100.47 618.275 ;
      RECT 100.755 0.17 101.525 0.43 ;
      RECT 101.265 0.17 101.525 8.7 ;
      RECT 100.755 0.17 101.015 16.7 ;
      RECT 100.245 0.3 100.505 4.63 ;
      RECT 100.765 617.545 100.965 618.275 ;
      RECT 101.265 617.545 101.465 618.275 ;
      RECT 101.765 617.545 101.965 618.275 ;
      RECT 102.26 617.545 102.46 618.275 ;
      RECT 103.08 617.545 103.28 618.275 ;
      RECT 103.575 617.545 103.775 618.275 ;
      RECT 104.075 617.545 104.275 618.275 ;
      RECT 104.575 617.545 104.775 618.275 ;
      RECT 105.07 617.545 105.27 618.275 ;
      RECT 105.89 617.545 106.09 618.275 ;
      RECT 106.385 617.545 106.585 618.275 ;
      RECT 106.885 617.545 107.085 618.275 ;
      RECT 107.385 617.545 107.585 618.275 ;
      RECT 107.485 0.3 107.745 4.63 ;
      RECT 108.505 0.165 109.275 0.425 ;
      RECT 108.505 0.165 108.765 8.825 ;
      RECT 109.015 0.165 109.275 8.825 ;
      RECT 107.88 617.545 108.08 618.275 ;
      RECT 107.995 0.3 108.255 4.63 ;
      RECT 108.7 617.545 108.9 618.275 ;
      RECT 109.195 617.545 109.395 618.275 ;
      RECT 109.695 617.545 109.895 618.275 ;
      RECT 109.935 0.52 110.195 4.5 ;
      RECT 110.195 617.545 110.395 618.275 ;
      RECT 110.69 617.545 110.89 618.275 ;
      RECT 111.51 617.545 111.71 618.275 ;
      RECT 112.005 617.545 112.205 618.275 ;
      RECT 112.505 617.545 112.705 618.275 ;
      RECT 113.005 617.545 113.205 618.275 ;
      RECT 113.5 617.545 113.7 618.275 ;
      RECT 114.32 617.545 114.52 618.275 ;
      RECT 114.815 617.545 115.015 618.275 ;
      RECT 115.315 617.545 115.515 618.275 ;
      RECT 115.815 617.545 116.015 618.275 ;
      RECT 116.31 617.545 116.51 618.275 ;
      RECT 117.13 617.545 117.33 618.275 ;
      RECT 117.625 617.545 117.825 618.275 ;
      RECT 118.125 617.545 118.325 618.275 ;
      RECT 118.625 617.545 118.825 618.275 ;
      RECT 119.12 617.545 119.32 618.275 ;
      RECT 119.94 617.545 120.14 618.275 ;
      RECT 120.435 617.545 120.635 618.275 ;
      RECT 120.935 617.545 121.135 618.275 ;
      RECT 121.435 617.545 121.635 618.275 ;
      RECT 121.93 617.545 122.13 618.275 ;
      RECT 122.75 617.545 122.95 618.275 ;
      RECT 123.705 0.16 124.475 0.42 ;
      RECT 124.215 0.16 124.475 4.63 ;
      RECT 123.705 0.16 123.965 8.82 ;
      RECT 123.245 617.545 123.445 618.275 ;
      RECT 123.745 617.545 123.945 618.275 ;
      RECT 124.245 617.545 124.445 618.275 ;
      RECT 124.74 617.545 124.94 618.275 ;
      RECT 124.725 0.3 124.985 4.63 ;
      RECT 125.235 0.3 125.495 4.63 ;
      RECT 125.56 617.545 125.76 618.275 ;
      RECT 126.055 617.545 126.255 618.275 ;
      RECT 126.555 617.545 126.755 618.275 ;
      RECT 128.24 0.16 129.01 0.42 ;
      RECT 128.24 0.16 128.5 8.82 ;
      RECT 128.75 0.16 129.01 8.82 ;
      RECT 127.055 617.545 127.255 618.275 ;
      RECT 127.55 617.545 127.75 618.275 ;
      RECT 128.37 617.545 128.57 618.275 ;
      RECT 128.865 617.545 129.065 618.275 ;
      RECT 129.26 0.3 129.52 4.63 ;
      RECT 129.365 617.545 129.565 618.275 ;
      RECT 129.77 0.3 130.03 4.63 ;
      RECT 129.865 617.545 130.065 618.275 ;
      RECT 130.36 617.545 130.56 618.275 ;
      RECT 130.775 0.52 131.035 10.655 ;
      RECT 131.18 617.545 131.38 618.275 ;
      RECT 131.675 617.545 131.875 618.275 ;
      RECT 131.71 0.52 131.97 4.5 ;
      RECT 132.175 617.545 132.375 618.275 ;
      RECT 132.675 617.545 132.875 618.275 ;
      RECT 133.17 617.545 133.37 618.275 ;
      RECT 134.415 0.165 135.185 0.425 ;
      RECT 134.415 0.165 134.675 8.825 ;
      RECT 134.925 0.165 135.185 8.825 ;
      RECT 133.99 617.545 134.19 618.275 ;
      RECT 134.485 617.545 134.685 618.275 ;
      RECT 134.985 617.545 135.185 618.275 ;
      RECT 135.485 617.545 135.685 618.275 ;
      RECT 135.435 0.3 135.695 4.63 ;
      RECT 135.98 617.545 136.18 618.275 ;
      RECT 135.945 0.3 136.205 8.23 ;
      RECT 136.8 617.545 137 618.275 ;
      RECT 137.295 617.545 137.495 618.275 ;
      RECT 137.71 0.52 137.97 7.94 ;
      RECT 137.795 617.545 137.995 618.275 ;
      RECT 138.295 617.545 138.495 618.275 ;
      RECT 138.79 617.545 138.99 618.275 ;
      RECT 139.24 0.52 139.5 10.655 ;
      RECT 140.105 0.17 140.875 0.43 ;
      RECT 140.615 0.17 140.875 11.38 ;
      RECT 140.105 0.17 140.365 16.7 ;
      RECT 139.61 617.545 139.81 618.275 ;
      RECT 140.105 617.545 140.305 618.275 ;
      RECT 140.605 617.545 140.805 618.275 ;
      RECT 141.105 617.545 141.305 618.275 ;
      RECT 141.6 617.545 141.8 618.275 ;
      RECT 142.42 617.545 142.62 618.275 ;
      RECT 143.675 0.17 144.445 0.43 ;
      RECT 144.185 0.17 144.445 8.7 ;
      RECT 143.675 0.17 143.935 16.7 ;
      RECT 142.915 617.545 143.115 618.275 ;
      RECT 143.415 617.545 143.615 618.275 ;
      RECT 143.915 617.545 144.115 618.275 ;
      RECT 144.41 617.545 144.61 618.275 ;
      RECT 144.695 0.3 144.955 4.63 ;
      RECT 145.23 617.545 145.43 618.275 ;
      RECT 145.715 0.17 146.485 0.43 ;
      RECT 146.225 0.17 146.485 8.7 ;
      RECT 145.715 0.17 145.975 16.7 ;
      RECT 145.205 0.3 145.465 4.63 ;
      RECT 145.725 617.545 145.925 618.275 ;
      RECT 146.225 617.545 146.425 618.275 ;
      RECT 146.725 617.545 146.925 618.275 ;
      RECT 147.22 617.545 147.42 618.275 ;
      RECT 148.04 617.545 148.24 618.275 ;
      RECT 148.535 617.545 148.735 618.275 ;
      RECT 149.035 617.545 149.235 618.275 ;
      RECT 149.535 617.545 149.735 618.275 ;
      RECT 150.03 617.545 150.23 618.275 ;
      RECT 150.85 617.545 151.05 618.275 ;
      RECT 151.345 617.545 151.545 618.275 ;
      RECT 151.845 617.545 152.045 618.275 ;
      RECT 152.345 617.545 152.545 618.275 ;
      RECT 152.445 0.3 152.705 4.63 ;
      RECT 153.465 0.165 154.235 0.425 ;
      RECT 153.465 0.165 153.725 8.825 ;
      RECT 153.975 0.165 154.235 8.825 ;
      RECT 152.84 617.545 153.04 618.275 ;
      RECT 152.955 0.3 153.215 4.63 ;
      RECT 153.66 617.545 153.86 618.275 ;
      RECT 154.155 617.545 154.355 618.275 ;
      RECT 154.655 617.545 154.855 618.275 ;
      RECT 154.895 0.52 155.155 4.5 ;
      RECT 155.155 617.545 155.355 618.275 ;
      RECT 155.65 617.545 155.85 618.275 ;
      RECT 156.47 617.545 156.67 618.275 ;
      RECT 156.965 617.545 157.165 618.275 ;
      RECT 157.465 617.545 157.665 618.275 ;
      RECT 157.965 617.545 158.165 618.275 ;
      RECT 158.46 617.545 158.66 618.275 ;
      RECT 159.28 617.545 159.48 618.275 ;
      RECT 159.775 617.545 159.975 618.275 ;
      RECT 160.275 617.545 160.475 618.275 ;
      RECT 160.775 617.545 160.975 618.275 ;
      RECT 161.27 617.545 161.47 618.275 ;
      RECT 162.09 617.545 162.29 618.275 ;
      RECT 162.585 617.545 162.785 618.275 ;
      RECT 163.085 617.545 163.285 618.275 ;
      RECT 163.585 617.545 163.785 618.275 ;
      RECT 164.08 617.545 164.28 618.275 ;
      RECT 164.9 617.545 165.1 618.275 ;
      RECT 165.395 617.545 165.595 618.275 ;
      RECT 165.895 617.545 166.095 618.275 ;
      RECT 166.395 617.545 166.595 618.275 ;
      RECT 166.89 617.545 167.09 618.275 ;
      RECT 167.71 617.545 167.91 618.275 ;
      RECT 168.665 0.16 169.435 0.42 ;
      RECT 169.175 0.16 169.435 4.63 ;
      RECT 168.665 0.16 168.925 8.82 ;
      RECT 168.205 617.545 168.405 618.275 ;
      RECT 168.705 617.545 168.905 618.275 ;
      RECT 169.205 617.545 169.405 618.275 ;
      RECT 169.7 617.545 169.9 618.275 ;
      RECT 169.685 0.3 169.945 4.63 ;
      RECT 170.195 0.3 170.455 4.63 ;
      RECT 170.52 617.545 170.72 618.275 ;
      RECT 171.015 617.545 171.215 618.275 ;
      RECT 171.515 617.545 171.715 618.275 ;
      RECT 173.2 0.16 173.97 0.42 ;
      RECT 173.2 0.16 173.46 8.82 ;
      RECT 173.71 0.16 173.97 8.82 ;
      RECT 172.015 617.545 172.215 618.275 ;
      RECT 172.51 617.545 172.71 618.275 ;
      RECT 173.33 617.545 173.53 618.275 ;
      RECT 173.825 617.545 174.025 618.275 ;
      RECT 174.22 0.3 174.48 4.63 ;
      RECT 174.325 617.545 174.525 618.275 ;
      RECT 174.73 0.3 174.99 4.63 ;
      RECT 174.825 617.545 175.025 618.275 ;
      RECT 175.32 617.545 175.52 618.275 ;
      RECT 175.735 0.52 175.995 10.655 ;
      RECT 176.14 617.545 176.34 618.275 ;
      RECT 176.635 617.545 176.835 618.275 ;
      RECT 176.67 0.52 176.93 4.5 ;
      RECT 177.135 617.545 177.335 618.275 ;
      RECT 177.635 617.545 177.835 618.275 ;
      RECT 178.13 617.545 178.33 618.275 ;
      RECT 179.375 0.165 180.145 0.425 ;
      RECT 179.375 0.165 179.635 8.825 ;
      RECT 179.885 0.165 180.145 8.825 ;
      RECT 178.95 617.545 179.15 618.275 ;
      RECT 179.445 617.545 179.645 618.275 ;
      RECT 179.945 617.545 180.145 618.275 ;
      RECT 180.445 617.545 180.645 618.275 ;
      RECT 180.395 0.3 180.655 4.63 ;
      RECT 180.94 617.545 181.14 618.275 ;
      RECT 180.905 0.3 181.165 8.23 ;
      RECT 181.76 617.545 181.96 618.275 ;
      RECT 182.255 617.545 182.455 618.275 ;
      RECT 182.67 0.52 182.93 7.94 ;
      RECT 182.755 617.545 182.955 618.275 ;
      RECT 183.255 617.545 183.455 618.275 ;
      RECT 183.75 617.545 183.95 618.275 ;
      RECT 184.2 0.52 184.46 10.655 ;
      RECT 185.065 0.17 185.835 0.43 ;
      RECT 185.575 0.17 185.835 11.38 ;
      RECT 185.065 0.17 185.325 16.7 ;
      RECT 184.57 617.545 184.77 618.275 ;
      RECT 185.065 617.545 185.265 618.275 ;
      RECT 185.565 617.545 185.765 618.275 ;
      RECT 186.065 617.545 186.265 618.275 ;
      RECT 186.56 617.545 186.76 618.275 ;
      RECT 187.38 617.545 187.58 618.275 ;
      RECT 188.635 0.17 189.405 0.43 ;
      RECT 189.145 0.17 189.405 8.7 ;
      RECT 188.635 0.17 188.895 16.7 ;
      RECT 187.875 617.545 188.075 618.275 ;
      RECT 188.375 617.545 188.575 618.275 ;
      RECT 188.875 617.545 189.075 618.275 ;
      RECT 189.37 617.545 189.57 618.275 ;
      RECT 189.655 0.3 189.915 4.63 ;
      RECT 190.19 617.545 190.39 618.275 ;
      RECT 190.675 0.17 191.445 0.43 ;
      RECT 191.185 0.17 191.445 8.7 ;
      RECT 190.675 0.17 190.935 16.7 ;
      RECT 190.165 0.3 190.425 4.63 ;
      RECT 190.685 617.545 190.885 618.275 ;
      RECT 191.185 617.545 191.385 618.275 ;
      RECT 191.685 617.545 191.885 618.275 ;
      RECT 192.18 617.545 192.38 618.275 ;
      RECT 193 617.545 193.2 618.275 ;
      RECT 193.495 617.545 193.695 618.275 ;
      RECT 193.995 617.545 194.195 618.275 ;
      RECT 194.495 617.545 194.695 618.275 ;
      RECT 194.99 617.545 195.19 618.275 ;
      RECT 195.81 617.545 196.01 618.275 ;
      RECT 196.305 617.545 196.505 618.275 ;
      RECT 196.805 617.545 197.005 618.275 ;
      RECT 197.305 617.545 197.505 618.275 ;
      RECT 197.405 0.3 197.665 4.63 ;
      RECT 198.425 0.165 199.195 0.425 ;
      RECT 198.425 0.165 198.685 8.825 ;
      RECT 198.935 0.165 199.195 8.825 ;
      RECT 197.8 617.545 198 618.275 ;
      RECT 197.915 0.3 198.175 4.63 ;
      RECT 198.62 617.545 198.82 618.275 ;
      RECT 199.115 617.545 199.315 618.275 ;
      RECT 199.615 617.545 199.815 618.275 ;
      RECT 199.855 0.52 200.115 4.5 ;
      RECT 200.115 617.545 200.315 618.275 ;
      RECT 200.61 617.545 200.81 618.275 ;
      RECT 201.43 617.545 201.63 618.275 ;
      RECT 201.925 617.545 202.125 618.275 ;
      RECT 202.425 617.545 202.625 618.275 ;
      RECT 202.925 617.545 203.125 618.275 ;
      RECT 203.42 617.545 203.62 618.275 ;
      RECT 204.24 617.545 204.44 618.275 ;
      RECT 204.735 617.545 204.935 618.275 ;
      RECT 205.235 617.545 205.435 618.275 ;
      RECT 205.735 617.545 205.935 618.275 ;
      RECT 206.23 617.545 206.43 618.275 ;
      RECT 207.05 617.545 207.25 618.275 ;
      RECT 207.545 617.545 207.745 618.275 ;
      RECT 208.045 617.545 208.245 618.275 ;
      RECT 208.545 617.545 208.745 618.275 ;
      RECT 209.04 617.545 209.24 618.275 ;
      RECT 209.86 617.545 210.06 618.275 ;
      RECT 210.355 617.545 210.555 618.275 ;
      RECT 210.855 617.545 211.055 618.275 ;
      RECT 211.355 617.545 211.555 618.275 ;
      RECT 211.85 617.545 212.05 618.275 ;
      RECT 212.67 617.545 212.87 618.275 ;
      RECT 213.625 0.16 214.395 0.42 ;
      RECT 214.135 0.16 214.395 4.63 ;
      RECT 213.625 0.16 213.885 8.82 ;
      RECT 213.165 617.545 213.365 618.275 ;
      RECT 213.665 617.545 213.865 618.275 ;
      RECT 214.165 617.545 214.365 618.275 ;
      RECT 214.66 617.545 214.86 618.275 ;
      RECT 214.645 0.3 214.905 4.63 ;
      RECT 215.155 0.3 215.415 4.63 ;
      RECT 215.48 617.545 215.68 618.275 ;
      RECT 215.975 617.545 216.175 618.275 ;
      RECT 216.475 617.545 216.675 618.275 ;
      RECT 218.16 0.16 218.93 0.42 ;
      RECT 218.16 0.16 218.42 8.82 ;
      RECT 218.67 0.16 218.93 8.82 ;
      RECT 216.975 617.545 217.175 618.275 ;
      RECT 217.47 617.545 217.67 618.275 ;
      RECT 218.29 617.545 218.49 618.275 ;
      RECT 218.785 617.545 218.985 618.275 ;
      RECT 219.18 0.3 219.44 4.63 ;
      RECT 219.285 617.545 219.485 618.275 ;
      RECT 219.69 0.3 219.95 4.63 ;
      RECT 219.785 617.545 219.985 618.275 ;
      RECT 220.28 617.545 220.48 618.275 ;
      RECT 220.695 0.52 220.955 10.655 ;
      RECT 221.1 617.545 221.3 618.275 ;
      RECT 221.595 617.545 221.795 618.275 ;
      RECT 221.63 0.52 221.89 4.5 ;
      RECT 222.095 617.545 222.295 618.275 ;
      RECT 222.595 617.545 222.795 618.275 ;
      RECT 223.09 617.545 223.29 618.275 ;
      RECT 224.335 0.165 225.105 0.425 ;
      RECT 224.335 0.165 224.595 8.825 ;
      RECT 224.845 0.165 225.105 8.825 ;
      RECT 223.91 617.545 224.11 618.275 ;
      RECT 224.405 617.545 224.605 618.275 ;
      RECT 224.905 617.545 225.105 618.275 ;
      RECT 225.405 617.545 225.605 618.275 ;
      RECT 225.355 0.3 225.615 4.63 ;
      RECT 225.9 617.545 226.1 618.275 ;
      RECT 225.865 0.3 226.125 8.23 ;
      RECT 226.72 617.545 226.92 618.275 ;
      RECT 227.215 617.545 227.415 618.275 ;
      RECT 227.63 0.52 227.89 7.94 ;
      RECT 227.715 617.545 227.915 618.275 ;
      RECT 228.215 617.545 228.415 618.275 ;
      RECT 228.71 617.545 228.91 618.275 ;
      RECT 229.16 0.52 229.42 10.655 ;
      RECT 230.025 0.17 230.795 0.43 ;
      RECT 230.535 0.17 230.795 11.38 ;
      RECT 230.025 0.17 230.285 16.7 ;
      RECT 229.53 617.545 229.73 618.275 ;
      RECT 230.025 617.545 230.225 618.275 ;
      RECT 230.525 617.545 230.725 618.275 ;
      RECT 231.025 617.545 231.225 618.275 ;
      RECT 231.52 617.545 231.72 618.275 ;
      RECT 232.34 617.545 232.54 618.275 ;
      RECT 233.595 0.17 234.365 0.43 ;
      RECT 234.105 0.17 234.365 8.7 ;
      RECT 233.595 0.17 233.855 16.7 ;
      RECT 232.835 617.545 233.035 618.275 ;
      RECT 233.335 617.545 233.535 618.275 ;
      RECT 233.835 617.545 234.035 618.275 ;
      RECT 234.33 617.545 234.53 618.275 ;
      RECT 234.615 0.3 234.875 4.63 ;
      RECT 235.15 617.545 235.35 618.275 ;
      RECT 235.635 0.17 236.405 0.43 ;
      RECT 236.145 0.17 236.405 8.7 ;
      RECT 235.635 0.17 235.895 16.7 ;
      RECT 235.125 0.3 235.385 4.63 ;
      RECT 235.645 617.545 235.845 618.275 ;
      RECT 236.145 617.545 236.345 618.275 ;
      RECT 236.645 617.545 236.845 618.275 ;
      RECT 237.14 617.545 237.34 618.275 ;
      RECT 237.96 617.545 238.16 618.275 ;
      RECT 238.455 617.545 238.655 618.275 ;
      RECT 238.955 617.545 239.155 618.275 ;
      RECT 239.455 617.545 239.655 618.275 ;
      RECT 239.95 617.545 240.15 618.275 ;
      RECT 240.77 617.545 240.97 618.275 ;
      RECT 241.265 617.545 241.465 618.275 ;
      RECT 241.765 617.545 241.965 618.275 ;
      RECT 242.265 617.545 242.465 618.275 ;
      RECT 242.365 0.3 242.625 4.63 ;
      RECT 243.385 0.165 244.155 0.425 ;
      RECT 243.385 0.165 243.645 8.825 ;
      RECT 243.895 0.165 244.155 8.825 ;
      RECT 242.76 617.545 242.96 618.275 ;
      RECT 242.875 0.3 243.135 4.63 ;
      RECT 243.58 617.545 243.78 618.275 ;
      RECT 244.075 617.545 244.275 618.275 ;
      RECT 244.575 617.545 244.775 618.275 ;
      RECT 244.815 0.52 245.075 4.5 ;
      RECT 245.075 617.545 245.275 618.275 ;
      RECT 245.57 617.545 245.77 618.275 ;
      RECT 246.39 617.545 246.59 618.275 ;
      RECT 246.885 617.545 247.085 618.275 ;
      RECT 247.385 617.545 247.585 618.275 ;
      RECT 247.885 617.545 248.085 618.275 ;
      RECT 248.38 617.545 248.58 618.275 ;
      RECT 249.2 617.545 249.4 618.275 ;
      RECT 249.695 617.545 249.895 618.275 ;
      RECT 250.195 617.545 250.395 618.275 ;
      RECT 250.695 617.545 250.895 618.275 ;
      RECT 251.19 617.545 251.39 618.275 ;
      RECT 252.01 617.545 252.21 618.275 ;
      RECT 252.505 617.545 252.705 618.275 ;
      RECT 253.005 617.545 253.205 618.275 ;
      RECT 253.505 617.545 253.705 618.275 ;
      RECT 254 617.545 254.2 618.275 ;
      RECT 254.82 617.545 255.02 618.275 ;
      RECT 255.315 617.545 255.515 618.275 ;
      RECT 255.815 617.545 256.015 618.275 ;
      RECT 256.315 617.545 256.515 618.275 ;
      RECT 256.81 617.545 257.01 618.275 ;
      RECT 257.63 617.545 257.83 618.275 ;
      RECT 258.585 0.16 259.355 0.42 ;
      RECT 259.095 0.16 259.355 4.63 ;
      RECT 258.585 0.16 258.845 8.82 ;
      RECT 258.125 617.545 258.325 618.275 ;
      RECT 258.625 617.545 258.825 618.275 ;
      RECT 259.125 617.545 259.325 618.275 ;
      RECT 259.62 617.545 259.82 618.275 ;
      RECT 259.605 0.3 259.865 4.63 ;
      RECT 260.115 0.3 260.375 4.63 ;
      RECT 260.44 617.545 260.64 618.275 ;
      RECT 260.935 617.545 261.135 618.275 ;
      RECT 261.435 617.545 261.635 618.275 ;
      RECT 263.12 0.16 263.89 0.42 ;
      RECT 263.12 0.16 263.38 8.82 ;
      RECT 263.63 0.16 263.89 8.82 ;
      RECT 261.935 617.545 262.135 618.275 ;
      RECT 262.43 617.545 262.63 618.275 ;
      RECT 263.25 617.545 263.45 618.275 ;
      RECT 263.745 617.545 263.945 618.275 ;
      RECT 264.14 0.3 264.4 4.63 ;
      RECT 264.245 617.545 264.445 618.275 ;
      RECT 264.65 0.3 264.91 4.63 ;
      RECT 264.745 617.545 264.945 618.275 ;
      RECT 265.24 617.545 265.44 618.275 ;
      RECT 265.655 0.52 265.915 10.655 ;
      RECT 266.06 617.545 266.26 618.275 ;
      RECT 266.555 617.545 266.755 618.275 ;
      RECT 266.59 0.52 266.85 4.5 ;
      RECT 267.055 617.545 267.255 618.275 ;
      RECT 267.555 617.545 267.755 618.275 ;
      RECT 268.05 617.545 268.25 618.275 ;
      RECT 269.295 0.165 270.065 0.425 ;
      RECT 269.295 0.165 269.555 8.825 ;
      RECT 269.805 0.165 270.065 8.825 ;
      RECT 268.87 617.545 269.07 618.275 ;
      RECT 269.365 617.545 269.565 618.275 ;
      RECT 269.865 617.545 270.065 618.275 ;
      RECT 270.365 617.545 270.565 618.275 ;
      RECT 270.315 0.3 270.575 4.63 ;
      RECT 270.86 617.545 271.06 618.275 ;
      RECT 270.825 0.3 271.085 8.23 ;
      RECT 271.68 617.545 271.88 618.275 ;
      RECT 272.175 617.545 272.375 618.275 ;
      RECT 272.59 0.52 272.85 7.94 ;
      RECT 272.675 617.545 272.875 618.275 ;
      RECT 273.175 617.545 273.375 618.275 ;
      RECT 273.67 617.545 273.87 618.275 ;
      RECT 274.12 0.52 274.38 10.655 ;
      RECT 274.985 0.17 275.755 0.43 ;
      RECT 275.495 0.17 275.755 11.38 ;
      RECT 274.985 0.17 275.245 16.7 ;
      RECT 274.49 617.545 274.69 618.275 ;
      RECT 274.985 617.545 275.185 618.275 ;
      RECT 275.485 617.545 275.685 618.275 ;
      RECT 275.985 617.545 276.185 618.275 ;
      RECT 276.48 617.545 276.68 618.275 ;
      RECT 277.3 617.545 277.5 618.275 ;
      RECT 278.555 0.17 279.325 0.43 ;
      RECT 279.065 0.17 279.325 8.7 ;
      RECT 278.555 0.17 278.815 16.7 ;
      RECT 277.795 617.545 277.995 618.275 ;
      RECT 278.295 617.545 278.495 618.275 ;
      RECT 278.795 617.545 278.995 618.275 ;
      RECT 279.29 617.545 279.49 618.275 ;
      RECT 279.575 0.3 279.835 4.63 ;
      RECT 280.11 617.545 280.31 618.275 ;
      RECT 280.595 0.17 281.365 0.43 ;
      RECT 281.105 0.17 281.365 8.7 ;
      RECT 280.595 0.17 280.855 16.7 ;
      RECT 280.085 0.3 280.345 4.63 ;
      RECT 280.605 617.545 280.805 618.275 ;
      RECT 281.105 617.545 281.305 618.275 ;
      RECT 281.605 617.545 281.805 618.275 ;
      RECT 282.1 617.545 282.3 618.275 ;
      RECT 282.92 617.545 283.12 618.275 ;
      RECT 283.415 617.545 283.615 618.275 ;
      RECT 283.915 617.545 284.115 618.275 ;
      RECT 284.415 617.545 284.615 618.275 ;
      RECT 284.91 617.545 285.11 618.275 ;
      RECT 285.73 617.545 285.93 618.275 ;
      RECT 286.225 617.545 286.425 618.275 ;
      RECT 286.725 617.545 286.925 618.275 ;
      RECT 287.225 617.545 287.425 618.275 ;
      RECT 287.325 0.3 287.585 4.63 ;
      RECT 288.345 0.165 289.115 0.425 ;
      RECT 288.345 0.165 288.605 8.825 ;
      RECT 288.855 0.165 289.115 8.825 ;
      RECT 287.72 617.545 287.92 618.275 ;
      RECT 287.835 0.3 288.095 4.63 ;
      RECT 288.54 617.545 288.74 618.275 ;
      RECT 289.035 617.545 289.235 618.275 ;
      RECT 289.535 617.545 289.735 618.275 ;
      RECT 289.775 0.52 290.035 4.5 ;
      RECT 290.035 617.545 290.235 618.275 ;
      RECT 290.53 617.545 290.73 618.275 ;
      RECT 291.35 617.545 291.55 618.275 ;
      RECT 291.845 617.545 292.045 618.275 ;
      RECT 292.345 617.545 292.545 618.275 ;
      RECT 292.845 617.545 293.045 618.275 ;
      RECT 293.34 617.545 293.54 618.275 ;
      RECT 294.16 617.545 294.36 618.275 ;
      RECT 294.655 617.545 294.855 618.275 ;
      RECT 295.155 617.545 295.355 618.275 ;
      RECT 295.655 617.545 295.855 618.275 ;
      RECT 296.15 617.545 296.35 618.275 ;
      RECT 296.97 617.545 297.17 618.275 ;
      RECT 297.465 617.545 297.665 618.275 ;
      RECT 297.965 617.545 298.165 618.275 ;
      RECT 298.465 617.545 298.665 618.275 ;
      RECT 298.96 617.545 299.16 618.275 ;
      RECT 299.78 617.545 299.98 618.275 ;
      RECT 300.275 617.545 300.475 618.275 ;
      RECT 300.775 617.545 300.975 618.275 ;
      RECT 301.275 617.545 301.475 618.275 ;
      RECT 301.77 617.545 301.97 618.275 ;
      RECT 302.59 617.545 302.79 618.275 ;
      RECT 303.545 0.16 304.315 0.42 ;
      RECT 304.055 0.16 304.315 4.63 ;
      RECT 303.545 0.16 303.805 8.82 ;
      RECT 303.085 617.545 303.285 618.275 ;
      RECT 303.585 617.545 303.785 618.275 ;
      RECT 304.085 617.545 304.285 618.275 ;
      RECT 304.58 617.545 304.78 618.275 ;
      RECT 304.565 0.3 304.825 4.63 ;
      RECT 305.075 0.3 305.335 4.63 ;
      RECT 305.4 617.545 305.6 618.275 ;
      RECT 305.895 617.545 306.095 618.275 ;
      RECT 306.395 617.545 306.595 618.275 ;
      RECT 308.08 0.16 308.85 0.42 ;
      RECT 308.08 0.16 308.34 8.82 ;
      RECT 308.59 0.16 308.85 8.82 ;
      RECT 306.895 617.545 307.095 618.275 ;
      RECT 307.39 617.545 307.59 618.275 ;
      RECT 308.21 617.545 308.41 618.275 ;
      RECT 308.705 617.545 308.905 618.275 ;
      RECT 309.1 0.3 309.36 4.63 ;
      RECT 309.205 617.545 309.405 618.275 ;
      RECT 309.61 0.3 309.87 4.63 ;
      RECT 309.705 617.545 309.905 618.275 ;
      RECT 310.2 617.545 310.4 618.275 ;
      RECT 310.615 0.52 310.875 10.655 ;
      RECT 311.02 617.545 311.22 618.275 ;
      RECT 311.515 617.545 311.715 618.275 ;
      RECT 311.55 0.52 311.81 4.5 ;
      RECT 312.015 617.545 312.215 618.275 ;
      RECT 312.515 617.545 312.715 618.275 ;
      RECT 313.01 617.545 313.21 618.275 ;
      RECT 314.255 0.165 315.025 0.425 ;
      RECT 314.255 0.165 314.515 8.825 ;
      RECT 314.765 0.165 315.025 8.825 ;
      RECT 313.83 617.545 314.03 618.275 ;
      RECT 314.325 617.545 314.525 618.275 ;
      RECT 314.825 617.545 315.025 618.275 ;
      RECT 315.325 617.545 315.525 618.275 ;
      RECT 315.275 0.3 315.535 4.63 ;
      RECT 315.82 617.545 316.02 618.275 ;
      RECT 315.785 0.3 316.045 8.23 ;
      RECT 316.64 617.545 316.84 618.275 ;
      RECT 317.135 617.545 317.335 618.275 ;
      RECT 317.55 0.52 317.81 7.94 ;
      RECT 317.635 617.545 317.835 618.275 ;
      RECT 318.135 617.545 318.335 618.275 ;
      RECT 318.63 617.545 318.83 618.275 ;
      RECT 319.08 0.52 319.34 10.655 ;
      RECT 319.945 0.17 320.715 0.43 ;
      RECT 320.455 0.17 320.715 11.38 ;
      RECT 319.945 0.17 320.205 16.7 ;
      RECT 319.45 617.545 319.65 618.275 ;
      RECT 319.945 617.545 320.145 618.275 ;
      RECT 320.445 617.545 320.645 618.275 ;
      RECT 320.945 617.545 321.145 618.275 ;
      RECT 321.44 617.545 321.64 618.275 ;
      RECT 322.26 617.545 322.46 618.275 ;
      RECT 323.515 0.17 324.285 0.43 ;
      RECT 324.025 0.17 324.285 8.7 ;
      RECT 323.515 0.17 323.775 16.7 ;
      RECT 322.755 617.545 322.955 618.275 ;
      RECT 323.255 617.545 323.455 618.275 ;
      RECT 323.755 617.545 323.955 618.275 ;
      RECT 324.25 617.545 324.45 618.275 ;
      RECT 324.535 0.3 324.795 4.63 ;
      RECT 325.07 617.545 325.27 618.275 ;
      RECT 325.555 0.17 326.325 0.43 ;
      RECT 326.065 0.17 326.325 8.7 ;
      RECT 325.555 0.17 325.815 16.7 ;
      RECT 325.045 0.3 325.305 4.63 ;
      RECT 325.565 617.545 325.765 618.275 ;
      RECT 326.065 617.545 326.265 618.275 ;
      RECT 326.565 617.545 326.765 618.275 ;
      RECT 327.06 617.545 327.26 618.275 ;
      RECT 327.88 617.545 328.08 618.275 ;
      RECT 328.375 617.545 328.575 618.275 ;
      RECT 328.875 617.545 329.075 618.275 ;
      RECT 329.375 617.545 329.575 618.275 ;
      RECT 329.87 617.545 330.07 618.275 ;
      RECT 330.69 617.545 330.89 618.275 ;
      RECT 331.185 617.545 331.385 618.275 ;
      RECT 331.685 617.545 331.885 618.275 ;
      RECT 332.185 617.545 332.385 618.275 ;
      RECT 332.285 0.3 332.545 4.63 ;
      RECT 333.305 0.165 334.075 0.425 ;
      RECT 333.305 0.165 333.565 8.825 ;
      RECT 333.815 0.165 334.075 8.825 ;
      RECT 332.68 617.545 332.88 618.275 ;
      RECT 332.795 0.3 333.055 4.63 ;
      RECT 333.5 617.545 333.7 618.275 ;
      RECT 333.995 617.545 334.195 618.275 ;
      RECT 334.495 617.545 334.695 618.275 ;
      RECT 334.735 0.52 334.995 4.5 ;
      RECT 334.995 617.545 335.195 618.275 ;
      RECT 335.49 617.545 335.69 618.275 ;
      RECT 336.31 617.545 336.51 618.275 ;
      RECT 336.805 617.545 337.005 618.275 ;
      RECT 337.305 617.545 337.505 618.275 ;
      RECT 337.805 617.545 338.005 618.275 ;
      RECT 338.3 617.545 338.5 618.275 ;
      RECT 339.12 617.545 339.32 618.275 ;
      RECT 339.615 617.545 339.815 618.275 ;
      RECT 340.115 617.545 340.315 618.275 ;
      RECT 340.615 617.545 340.815 618.275 ;
      RECT 341.11 617.545 341.31 618.275 ;
      RECT 341.93 617.545 342.13 618.275 ;
      RECT 342.425 617.545 342.625 618.275 ;
      RECT 342.925 617.545 343.125 618.275 ;
      RECT 343.425 617.545 343.625 618.275 ;
      RECT 343.92 617.545 344.12 618.275 ;
      RECT 344.74 617.545 344.94 618.275 ;
      RECT 345.235 617.545 345.435 618.275 ;
      RECT 345.735 617.545 345.935 618.275 ;
      RECT 346.235 617.545 346.435 618.275 ;
      RECT 346.73 617.545 346.93 618.275 ;
      RECT 347.55 617.545 347.75 618.275 ;
      RECT 348.505 0.16 349.275 0.42 ;
      RECT 349.015 0.16 349.275 4.63 ;
      RECT 348.505 0.16 348.765 8.82 ;
      RECT 348.045 617.545 348.245 618.275 ;
      RECT 348.545 617.545 348.745 618.275 ;
      RECT 349.045 617.545 349.245 618.275 ;
      RECT 349.54 617.545 349.74 618.275 ;
      RECT 349.525 0.3 349.785 4.63 ;
      RECT 350.035 0.3 350.295 4.63 ;
      RECT 350.36 617.545 350.56 618.275 ;
      RECT 350.855 617.545 351.055 618.275 ;
      RECT 351.355 617.545 351.555 618.275 ;
      RECT 353.04 0.16 353.81 0.42 ;
      RECT 353.04 0.16 353.3 8.82 ;
      RECT 353.55 0.16 353.81 8.82 ;
      RECT 351.855 617.545 352.055 618.275 ;
      RECT 352.35 617.545 352.55 618.275 ;
      RECT 353.17 617.545 353.37 618.275 ;
      RECT 353.665 617.545 353.865 618.275 ;
      RECT 354.06 0.3 354.32 4.63 ;
      RECT 354.165 617.545 354.365 618.275 ;
      RECT 354.57 0.3 354.83 4.63 ;
      RECT 354.665 617.545 354.865 618.275 ;
      RECT 355.16 617.545 355.36 618.275 ;
      RECT 355.575 0.52 355.835 10.655 ;
      RECT 355.98 617.545 356.18 618.275 ;
      RECT 356.475 617.545 356.675 618.275 ;
      RECT 356.51 0.52 356.77 4.5 ;
      RECT 356.975 617.545 357.175 618.275 ;
      RECT 357.475 617.545 357.675 618.275 ;
      RECT 357.97 617.545 358.17 618.275 ;
      RECT 359.215 0.165 359.985 0.425 ;
      RECT 359.215 0.165 359.475 8.825 ;
      RECT 359.725 0.165 359.985 8.825 ;
      RECT 358.79 617.545 358.99 618.275 ;
      RECT 359.285 617.545 359.485 618.275 ;
      RECT 359.785 617.545 359.985 618.275 ;
      RECT 360.285 617.545 360.485 618.275 ;
      RECT 360.235 0.3 360.495 4.63 ;
      RECT 360.78 617.545 360.98 618.275 ;
      RECT 360.745 0.3 361.005 8.23 ;
      RECT 361.6 617.545 361.8 618.275 ;
      RECT 362.095 617.545 362.295 618.275 ;
      RECT 362.51 0.52 362.77 7.94 ;
      RECT 362.595 617.545 362.795 618.275 ;
      RECT 363.095 617.545 363.295 618.275 ;
      RECT 363.59 617.545 363.79 618.275 ;
      RECT 364.04 0.52 364.3 10.655 ;
      RECT 364.905 0.17 365.675 0.43 ;
      RECT 365.415 0.17 365.675 11.38 ;
      RECT 364.905 0.17 365.165 16.7 ;
      RECT 364.41 617.545 364.61 618.275 ;
      RECT 364.905 617.545 365.105 618.275 ;
      RECT 365.405 617.545 365.605 618.275 ;
      RECT 365.905 617.545 366.105 618.275 ;
      RECT 366.4 617.545 366.6 618.275 ;
      RECT 367.22 617.545 367.42 618.275 ;
      RECT 368.475 0.17 369.245 0.43 ;
      RECT 368.985 0.17 369.245 8.7 ;
      RECT 368.475 0.17 368.735 16.7 ;
      RECT 367.715 617.545 367.915 618.275 ;
      RECT 368.215 617.545 368.415 618.275 ;
      RECT 368.715 617.545 368.915 618.275 ;
      RECT 369.21 617.545 369.41 618.275 ;
      RECT 369.495 0.3 369.755 4.63 ;
      RECT 370.03 617.545 370.23 618.275 ;
      RECT 370.515 0.17 371.285 0.43 ;
      RECT 371.025 0.17 371.285 8.7 ;
      RECT 370.515 0.17 370.775 16.7 ;
      RECT 370.005 0.3 370.265 4.63 ;
      RECT 370.525 617.545 370.725 618.275 ;
      RECT 371.025 617.545 371.225 618.275 ;
      RECT 371.525 617.545 371.725 618.275 ;
      RECT 372.02 617.545 372.22 618.275 ;
      RECT 372.84 617.545 373.04 618.275 ;
      RECT 373.335 617.545 373.535 618.275 ;
      RECT 373.835 617.545 374.035 618.275 ;
      RECT 374.335 617.545 374.535 618.275 ;
      RECT 374.83 617.545 375.03 618.275 ;
      RECT 375.65 617.545 375.85 618.275 ;
      RECT 376.145 617.545 376.345 618.275 ;
      RECT 376.645 617.545 376.845 618.275 ;
      RECT 377.145 617.545 377.345 618.275 ;
      RECT 377.245 0.3 377.505 4.63 ;
      RECT 378.265 0.165 379.035 0.425 ;
      RECT 378.265 0.165 378.525 8.825 ;
      RECT 378.775 0.165 379.035 8.825 ;
      RECT 377.64 617.545 377.84 618.275 ;
      RECT 377.755 0.3 378.015 4.63 ;
      RECT 378.46 617.545 378.66 618.275 ;
      RECT 378.955 617.545 379.155 618.275 ;
      RECT 379.455 617.545 379.655 618.275 ;
      RECT 379.695 0.52 379.955 4.5 ;
      RECT 379.955 617.545 380.155 618.275 ;
      RECT 380.45 617.545 380.65 618.275 ;
      RECT 381.27 617.545 381.47 618.275 ;
      RECT 381.765 617.545 381.965 618.275 ;
      RECT 382.265 617.545 382.465 618.275 ;
      RECT 382.765 617.545 382.965 618.275 ;
      RECT 383.26 617.545 383.46 618.275 ;
      RECT 384.08 617.545 384.28 618.275 ;
      RECT 384.575 617.545 384.775 618.275 ;
      RECT 385.075 617.545 385.275 618.275 ;
      RECT 385.575 617.545 385.775 618.275 ;
      RECT 386.07 617.545 386.27 618.275 ;
      RECT 386.89 617.545 387.09 618.275 ;
      RECT 387.385 617.545 387.585 618.275 ;
      RECT 387.885 617.545 388.085 618.275 ;
      RECT 388.385 617.545 388.585 618.275 ;
      RECT 388.88 617.545 389.08 618.275 ;
      RECT 389.7 617.545 389.9 618.275 ;
      RECT 390.195 617.545 390.395 618.275 ;
      RECT 390.695 617.545 390.895 618.275 ;
      RECT 391.195 617.545 391.395 618.275 ;
      RECT 391.69 617.545 391.89 618.275 ;
      RECT 392.51 617.545 392.71 618.275 ;
      RECT 393.465 0.16 394.235 0.42 ;
      RECT 393.975 0.16 394.235 4.63 ;
      RECT 393.465 0.16 393.725 8.82 ;
      RECT 393.005 617.545 393.205 618.275 ;
      RECT 393.505 617.545 393.705 618.275 ;
      RECT 394.005 617.545 394.205 618.275 ;
      RECT 394.5 617.545 394.7 618.275 ;
      RECT 394.485 0.3 394.745 4.63 ;
      RECT 394.995 0.3 395.255 4.63 ;
      RECT 395.32 617.545 395.52 618.275 ;
      RECT 395.815 617.545 396.015 618.275 ;
      RECT 396.315 617.545 396.515 618.275 ;
      RECT 398 0.16 398.77 0.42 ;
      RECT 398 0.16 398.26 8.82 ;
      RECT 398.51 0.16 398.77 8.82 ;
      RECT 396.815 617.545 397.015 618.275 ;
      RECT 397.31 617.545 397.51 618.275 ;
      RECT 398.13 617.545 398.33 618.275 ;
      RECT 398.625 617.545 398.825 618.275 ;
      RECT 399.02 0.3 399.28 4.63 ;
      RECT 399.125 617.545 399.325 618.275 ;
      RECT 399.53 0.3 399.79 4.63 ;
      RECT 399.625 617.545 399.825 618.275 ;
      RECT 400.12 617.545 400.32 618.275 ;
      RECT 400.535 0.52 400.795 10.655 ;
      RECT 400.94 617.545 401.14 618.275 ;
      RECT 401.435 617.545 401.635 618.275 ;
      RECT 401.47 0.52 401.73 4.5 ;
      RECT 401.935 617.545 402.135 618.275 ;
      RECT 402.435 617.545 402.635 618.275 ;
      RECT 402.93 617.545 403.13 618.275 ;
      RECT 404.175 0.165 404.945 0.425 ;
      RECT 404.175 0.165 404.435 8.825 ;
      RECT 404.685 0.165 404.945 8.825 ;
      RECT 403.75 617.545 403.95 618.275 ;
      RECT 404.245 617.545 404.445 618.275 ;
      RECT 404.745 617.545 404.945 618.275 ;
      RECT 405.245 617.545 405.445 618.275 ;
      RECT 405.195 0.3 405.455 4.63 ;
      RECT 405.74 617.545 405.94 618.275 ;
      RECT 405.705 0.3 405.965 8.23 ;
      RECT 406.56 617.545 406.76 618.275 ;
      RECT 407.055 617.545 407.255 618.275 ;
      RECT 407.47 0.52 407.73 7.94 ;
      RECT 407.555 617.545 407.755 618.275 ;
      RECT 408.055 617.545 408.255 618.275 ;
      RECT 408.55 617.545 408.75 618.275 ;
      RECT 409 0.52 409.26 10.655 ;
      RECT 409.865 0.17 410.635 0.43 ;
      RECT 410.375 0.17 410.635 11.38 ;
      RECT 409.865 0.17 410.125 16.7 ;
      RECT 409.37 617.545 409.57 618.275 ;
      RECT 409.865 617.545 410.065 618.275 ;
      RECT 410.365 617.545 410.565 618.275 ;
      RECT 410.865 617.545 411.065 618.275 ;
      RECT 411.36 617.545 411.56 618.275 ;
      RECT 412.18 617.545 412.38 618.275 ;
      RECT 413.435 0.17 414.205 0.43 ;
      RECT 413.945 0.17 414.205 8.7 ;
      RECT 413.435 0.17 413.695 16.7 ;
      RECT 412.675 617.545 412.875 618.275 ;
      RECT 413.175 617.545 413.375 618.275 ;
      RECT 413.675 617.545 413.875 618.275 ;
      RECT 414.17 617.545 414.37 618.275 ;
      RECT 414.455 0.3 414.715 4.63 ;
      RECT 414.99 617.545 415.19 618.275 ;
      RECT 415.475 0.17 416.245 0.43 ;
      RECT 415.985 0.17 416.245 8.7 ;
      RECT 415.475 0.17 415.735 16.7 ;
      RECT 414.965 0.3 415.225 4.63 ;
      RECT 415.485 617.545 415.685 618.275 ;
      RECT 415.985 617.545 416.185 618.275 ;
      RECT 416.485 617.545 416.685 618.275 ;
      RECT 416.98 617.545 417.18 618.275 ;
      RECT 417.8 617.545 418 618.275 ;
      RECT 418.295 617.545 418.495 618.275 ;
      RECT 418.795 617.545 418.995 618.275 ;
      RECT 419.295 617.545 419.495 618.275 ;
      RECT 419.79 617.545 419.99 618.275 ;
      RECT 420.61 617.545 420.81 618.275 ;
      RECT 421.105 617.545 421.305 618.275 ;
      RECT 421.605 617.545 421.805 618.275 ;
      RECT 422.105 617.545 422.305 618.275 ;
      RECT 422.205 0.3 422.465 4.63 ;
      RECT 423.225 0.165 423.995 0.425 ;
      RECT 423.225 0.165 423.485 8.825 ;
      RECT 423.735 0.165 423.995 8.825 ;
      RECT 422.6 617.545 422.8 618.275 ;
      RECT 422.715 0.3 422.975 4.63 ;
      RECT 423.42 617.545 423.62 618.275 ;
      RECT 423.915 617.545 424.115 618.275 ;
      RECT 424.415 617.545 424.615 618.275 ;
      RECT 424.655 0.52 424.915 4.5 ;
      RECT 424.915 617.545 425.115 618.275 ;
      RECT 425.41 617.545 425.61 618.275 ;
      RECT 426.23 617.545 426.43 618.275 ;
      RECT 426.725 617.545 426.925 618.275 ;
      RECT 427.225 617.545 427.425 618.275 ;
      RECT 427.725 617.545 427.925 618.275 ;
      RECT 428.22 617.545 428.42 618.275 ;
      RECT 429.04 617.545 429.24 618.275 ;
      RECT 429.535 617.545 429.735 618.275 ;
      RECT 430.035 617.545 430.235 618.275 ;
      RECT 430.535 617.545 430.735 618.275 ;
      RECT 431.03 617.545 431.23 618.275 ;
      RECT 431.85 617.545 432.05 618.275 ;
      RECT 432.345 617.545 432.545 618.275 ;
      RECT 432.845 617.545 433.045 618.275 ;
      RECT 433.345 617.545 433.545 618.275 ;
      RECT 433.84 617.545 434.04 618.275 ;
      RECT 434.66 617.545 434.86 618.275 ;
      RECT 435.155 617.545 435.355 618.275 ;
      RECT 435.655 617.545 435.855 618.275 ;
      RECT 436.155 617.545 436.355 618.275 ;
      RECT 436.65 617.545 436.85 618.275 ;
      RECT 437.47 617.545 437.67 618.275 ;
      RECT 438.425 0.16 439.195 0.42 ;
      RECT 438.935 0.16 439.195 4.63 ;
      RECT 438.425 0.16 438.685 8.82 ;
      RECT 437.965 617.545 438.165 618.275 ;
      RECT 438.465 617.545 438.665 618.275 ;
      RECT 438.965 617.545 439.165 618.275 ;
      RECT 439.46 617.545 439.66 618.275 ;
      RECT 439.445 0.3 439.705 4.63 ;
      RECT 439.955 0.3 440.215 4.63 ;
      RECT 440.28 617.545 440.48 618.275 ;
      RECT 440.775 617.545 440.975 618.275 ;
      RECT 441.275 617.545 441.475 618.275 ;
      RECT 442.96 0.16 443.73 0.42 ;
      RECT 442.96 0.16 443.22 8.82 ;
      RECT 443.47 0.16 443.73 8.82 ;
      RECT 441.775 617.545 441.975 618.275 ;
      RECT 442.27 617.545 442.47 618.275 ;
      RECT 443.09 617.545 443.29 618.275 ;
      RECT 443.585 617.545 443.785 618.275 ;
      RECT 443.98 0.3 444.24 4.63 ;
      RECT 444.085 617.545 444.285 618.275 ;
      RECT 444.49 0.3 444.75 4.63 ;
      RECT 444.585 617.545 444.785 618.275 ;
      RECT 445.08 617.545 445.28 618.275 ;
      RECT 445.495 0.52 445.755 10.655 ;
      RECT 445.9 617.545 446.1 618.275 ;
      RECT 446.395 617.545 446.595 618.275 ;
      RECT 446.43 0.52 446.69 4.5 ;
      RECT 446.895 617.545 447.095 618.275 ;
      RECT 447.395 617.545 447.595 618.275 ;
      RECT 447.89 617.545 448.09 618.275 ;
      RECT 449.135 0.165 449.905 0.425 ;
      RECT 449.135 0.165 449.395 8.825 ;
      RECT 449.645 0.165 449.905 8.825 ;
      RECT 448.71 617.545 448.91 618.275 ;
      RECT 449.205 617.545 449.405 618.275 ;
      RECT 449.705 617.545 449.905 618.275 ;
      RECT 450.205 617.545 450.405 618.275 ;
      RECT 450.155 0.3 450.415 4.63 ;
      RECT 450.7 617.545 450.9 618.275 ;
      RECT 450.665 0.3 450.925 8.23 ;
      RECT 451.52 617.545 451.72 618.275 ;
      RECT 452.015 617.545 452.215 618.275 ;
      RECT 452.43 0.52 452.69 7.94 ;
      RECT 452.515 617.545 452.715 618.275 ;
      RECT 453.015 617.545 453.215 618.275 ;
      RECT 453.51 617.545 453.71 618.275 ;
      RECT 453.96 0.52 454.22 10.655 ;
      RECT 454.825 0.17 455.595 0.43 ;
      RECT 455.335 0.17 455.595 11.38 ;
      RECT 454.825 0.17 455.085 16.7 ;
      RECT 454.33 617.545 454.53 618.275 ;
      RECT 454.825 617.545 455.025 618.275 ;
      RECT 455.325 617.545 455.525 618.275 ;
      RECT 455.825 617.545 456.025 618.275 ;
      RECT 456.32 617.545 456.52 618.275 ;
      RECT 457.14 617.545 457.34 618.275 ;
      RECT 458.395 0.17 459.165 0.43 ;
      RECT 458.905 0.17 459.165 8.7 ;
      RECT 458.395 0.17 458.655 16.7 ;
      RECT 457.635 617.545 457.835 618.275 ;
      RECT 458.135 617.545 458.335 618.275 ;
      RECT 458.635 617.545 458.835 618.275 ;
      RECT 459.13 617.545 459.33 618.275 ;
      RECT 459.415 0.3 459.675 4.63 ;
      RECT 459.95 617.545 460.15 618.275 ;
      RECT 460.435 0.17 461.205 0.43 ;
      RECT 460.945 0.17 461.205 8.7 ;
      RECT 460.435 0.17 460.695 16.7 ;
      RECT 459.925 0.3 460.185 4.63 ;
      RECT 460.445 617.545 460.645 618.275 ;
      RECT 460.945 617.545 461.145 618.275 ;
      RECT 461.445 617.545 461.645 618.275 ;
      RECT 461.94 617.545 462.14 618.275 ;
      RECT 462.76 617.545 462.96 618.275 ;
      RECT 463.255 617.545 463.455 618.275 ;
      RECT 463.755 617.545 463.955 618.275 ;
      RECT 464.255 617.545 464.455 618.275 ;
      RECT 464.75 617.545 464.95 618.275 ;
      RECT 465.57 617.545 465.77 618.275 ;
      RECT 466.065 617.545 466.265 618.275 ;
      RECT 466.565 617.545 466.765 618.275 ;
      RECT 467.065 617.545 467.265 618.275 ;
      RECT 467.165 0.3 467.425 4.63 ;
      RECT 468.185 0.165 468.955 0.425 ;
      RECT 468.185 0.165 468.445 8.825 ;
      RECT 468.695 0.165 468.955 8.825 ;
      RECT 467.56 617.545 467.76 618.275 ;
      RECT 467.675 0.3 467.935 4.63 ;
      RECT 468.38 617.545 468.58 618.275 ;
      RECT 468.875 617.545 469.075 618.275 ;
      RECT 469.375 617.545 469.575 618.275 ;
      RECT 469.615 0.52 469.875 4.5 ;
      RECT 469.875 617.545 470.075 618.275 ;
      RECT 470.37 617.545 470.57 618.275 ;
      RECT 471.19 617.545 471.39 618.275 ;
      RECT 471.685 617.545 471.885 618.275 ;
      RECT 472.185 617.545 472.385 618.275 ;
      RECT 472.685 617.545 472.885 618.275 ;
      RECT 473.18 617.545 473.38 618.275 ;
      RECT 474 617.545 474.2 618.275 ;
      RECT 474.495 617.545 474.695 618.275 ;
      RECT 474.995 617.545 475.195 618.275 ;
      RECT 475.495 617.545 475.695 618.275 ;
      RECT 475.99 617.545 476.19 618.275 ;
      RECT 476.81 617.545 477.01 618.275 ;
      RECT 477.305 617.545 477.505 618.275 ;
      RECT 477.805 617.545 478.005 618.275 ;
      RECT 478.305 617.545 478.505 618.275 ;
      RECT 478.8 617.545 479 618.275 ;
      RECT 479.62 617.545 479.82 618.275 ;
      RECT 480.115 617.545 480.315 618.275 ;
      RECT 480.615 617.545 480.815 618.275 ;
      RECT 481.115 617.545 481.315 618.275 ;
      RECT 481.61 617.545 481.81 618.275 ;
      RECT 482.43 617.545 482.63 618.275 ;
      RECT 483.385 0.16 484.155 0.42 ;
      RECT 483.895 0.16 484.155 4.63 ;
      RECT 483.385 0.16 483.645 8.82 ;
      RECT 482.925 617.545 483.125 618.275 ;
      RECT 483.425 617.545 483.625 618.275 ;
      RECT 483.925 617.545 484.125 618.275 ;
      RECT 484.42 617.545 484.62 618.275 ;
      RECT 484.405 0.3 484.665 4.63 ;
      RECT 484.915 0.3 485.175 4.63 ;
      RECT 485.24 617.545 485.44 618.275 ;
      RECT 485.735 617.545 485.935 618.275 ;
      RECT 486.235 617.545 486.435 618.275 ;
      RECT 487.92 0.16 488.69 0.42 ;
      RECT 487.92 0.16 488.18 8.82 ;
      RECT 488.43 0.16 488.69 8.82 ;
      RECT 486.735 617.545 486.935 618.275 ;
      RECT 487.23 617.545 487.43 618.275 ;
      RECT 488.05 617.545 488.25 618.275 ;
      RECT 488.545 617.545 488.745 618.275 ;
      RECT 488.94 0.3 489.2 4.63 ;
      RECT 489.045 617.545 489.245 618.275 ;
      RECT 489.45 0.3 489.71 4.63 ;
      RECT 489.545 617.545 489.745 618.275 ;
      RECT 490.04 617.545 490.24 618.275 ;
      RECT 490.455 0.52 490.715 10.655 ;
      RECT 490.86 617.545 491.06 618.275 ;
      RECT 491.355 617.545 491.555 618.275 ;
      RECT 491.39 0.52 491.65 4.5 ;
      RECT 491.855 617.545 492.055 618.275 ;
      RECT 492.355 617.545 492.555 618.275 ;
      RECT 492.85 617.545 493.05 618.275 ;
      RECT 494.095 0.165 494.865 0.425 ;
      RECT 494.095 0.165 494.355 8.825 ;
      RECT 494.605 0.165 494.865 8.825 ;
      RECT 493.67 617.545 493.87 618.275 ;
      RECT 494.165 617.545 494.365 618.275 ;
      RECT 494.665 617.545 494.865 618.275 ;
      RECT 495.165 617.545 495.365 618.275 ;
      RECT 495.115 0.3 495.375 4.63 ;
      RECT 495.66 617.545 495.86 618.275 ;
      RECT 495.625 0.3 495.885 8.23 ;
      RECT 496.48 617.545 496.68 618.275 ;
      RECT 496.975 617.545 497.175 618.275 ;
      RECT 497.39 0.52 497.65 7.94 ;
      RECT 497.475 617.545 497.675 618.275 ;
      RECT 497.975 617.545 498.175 618.275 ;
      RECT 498.47 617.545 498.67 618.275 ;
      RECT 498.92 0.52 499.18 10.655 ;
      RECT 499.785 0.17 500.555 0.43 ;
      RECT 500.295 0.17 500.555 11.38 ;
      RECT 499.785 0.17 500.045 16.7 ;
      RECT 499.29 617.545 499.49 618.275 ;
      RECT 499.785 617.545 499.985 618.275 ;
      RECT 500.285 617.545 500.485 618.275 ;
      RECT 500.785 617.545 500.985 618.275 ;
      RECT 501.28 617.545 501.48 618.275 ;
      RECT 502.1 617.545 502.3 618.275 ;
      RECT 503.355 0.17 504.125 0.43 ;
      RECT 503.865 0.17 504.125 8.7 ;
      RECT 503.355 0.17 503.615 16.7 ;
      RECT 502.595 617.545 502.795 618.275 ;
      RECT 503.095 617.545 503.295 618.275 ;
      RECT 503.595 617.545 503.795 618.275 ;
      RECT 504.09 617.545 504.29 618.275 ;
      RECT 504.375 0.3 504.635 4.63 ;
      RECT 504.91 617.545 505.11 618.275 ;
      RECT 505.395 0.17 506.165 0.43 ;
      RECT 505.905 0.17 506.165 8.7 ;
      RECT 505.395 0.17 505.655 16.7 ;
      RECT 504.885 0.3 505.145 4.63 ;
      RECT 505.405 617.545 505.605 618.275 ;
      RECT 505.905 617.545 506.105 618.275 ;
      RECT 506.405 617.545 506.605 618.275 ;
      RECT 506.9 617.545 507.1 618.275 ;
      RECT 507.72 617.545 507.92 618.275 ;
      RECT 508.215 617.545 508.415 618.275 ;
      RECT 508.715 617.545 508.915 618.275 ;
      RECT 509.215 617.545 509.415 618.275 ;
      RECT 509.71 617.545 509.91 618.275 ;
      RECT 510.53 617.545 510.73 618.275 ;
      RECT 511.025 617.545 511.225 618.275 ;
      RECT 511.525 617.545 511.725 618.275 ;
      RECT 512.025 617.545 512.225 618.275 ;
      RECT 512.125 0.3 512.385 4.63 ;
      RECT 513.145 0.165 513.915 0.425 ;
      RECT 513.145 0.165 513.405 8.825 ;
      RECT 513.655 0.165 513.915 8.825 ;
      RECT 512.52 617.545 512.72 618.275 ;
      RECT 512.635 0.3 512.895 4.63 ;
      RECT 513.34 617.545 513.54 618.275 ;
      RECT 513.835 617.545 514.035 618.275 ;
      RECT 514.335 617.545 514.535 618.275 ;
      RECT 514.575 0.52 514.835 4.5 ;
      RECT 514.835 617.545 515.035 618.275 ;
      RECT 515.33 617.545 515.53 618.275 ;
      RECT 516.15 617.545 516.35 618.275 ;
      RECT 516.645 617.545 516.845 618.275 ;
      RECT 517.145 617.545 517.345 618.275 ;
      RECT 517.645 617.545 517.845 618.275 ;
      RECT 518.14 617.545 518.34 618.275 ;
      RECT 518.96 617.545 519.16 618.275 ;
      RECT 519.455 617.545 519.655 618.275 ;
      RECT 519.955 617.545 520.155 618.275 ;
      RECT 520.455 617.545 520.655 618.275 ;
      RECT 520.95 617.545 521.15 618.275 ;
      RECT 521.77 617.545 521.97 618.275 ;
      RECT 522.265 617.545 522.465 618.275 ;
      RECT 522.765 617.545 522.965 618.275 ;
      RECT 523.265 617.545 523.465 618.275 ;
      RECT 523.76 617.545 523.96 618.275 ;
      RECT 524.58 617.545 524.78 618.275 ;
      RECT 525.075 617.545 525.275 618.275 ;
      RECT 525.575 617.545 525.775 618.275 ;
      RECT 526.075 617.545 526.275 618.275 ;
      RECT 526.57 617.545 526.77 618.275 ;
      RECT 527.39 617.545 527.59 618.275 ;
      RECT 528.345 0.16 529.115 0.42 ;
      RECT 528.855 0.16 529.115 4.63 ;
      RECT 528.345 0.16 528.605 8.82 ;
      RECT 527.885 617.545 528.085 618.275 ;
      RECT 528.385 617.545 528.585 618.275 ;
      RECT 528.885 617.545 529.085 618.275 ;
      RECT 529.38 617.545 529.58 618.275 ;
      RECT 529.365 0.3 529.625 4.63 ;
      RECT 529.875 0.3 530.135 4.63 ;
      RECT 530.2 617.545 530.4 618.275 ;
      RECT 530.695 617.545 530.895 618.275 ;
      RECT 531.195 617.545 531.395 618.275 ;
      RECT 532.88 0.16 533.65 0.42 ;
      RECT 532.88 0.16 533.14 8.82 ;
      RECT 533.39 0.16 533.65 8.82 ;
      RECT 531.695 617.545 531.895 618.275 ;
      RECT 532.19 617.545 532.39 618.275 ;
      RECT 533.01 617.545 533.21 618.275 ;
      RECT 533.505 617.545 533.705 618.275 ;
      RECT 533.9 0.3 534.16 4.63 ;
      RECT 534.005 617.545 534.205 618.275 ;
      RECT 534.41 0.3 534.67 4.63 ;
      RECT 534.505 617.545 534.705 618.275 ;
      RECT 535 617.545 535.2 618.275 ;
      RECT 535.415 0.52 535.675 10.655 ;
      RECT 535.82 617.545 536.02 618.275 ;
      RECT 536.315 617.545 536.515 618.275 ;
      RECT 536.35 0.52 536.61 4.5 ;
      RECT 536.815 617.545 537.015 618.275 ;
      RECT 537.315 617.545 537.515 618.275 ;
      RECT 537.81 617.545 538.01 618.275 ;
      RECT 539.055 0.165 539.825 0.425 ;
      RECT 539.055 0.165 539.315 8.825 ;
      RECT 539.565 0.165 539.825 8.825 ;
      RECT 538.63 617.545 538.83 618.275 ;
      RECT 539.125 617.545 539.325 618.275 ;
      RECT 539.625 617.545 539.825 618.275 ;
      RECT 540.125 617.545 540.325 618.275 ;
      RECT 540.075 0.3 540.335 4.63 ;
      RECT 540.62 617.545 540.82 618.275 ;
      RECT 540.585 0.3 540.845 8.23 ;
      RECT 541.44 617.545 541.64 618.275 ;
      RECT 541.935 617.545 542.135 618.275 ;
      RECT 542.35 0.52 542.61 7.94 ;
      RECT 542.435 617.545 542.635 618.275 ;
      RECT 542.935 617.545 543.135 618.275 ;
      RECT 543.43 617.545 543.63 618.275 ;
      RECT 543.88 0.52 544.14 10.655 ;
      RECT 544.745 0.17 545.515 0.43 ;
      RECT 545.255 0.17 545.515 11.38 ;
      RECT 544.745 0.17 545.005 16.7 ;
      RECT 544.25 617.545 544.45 618.275 ;
      RECT 544.745 617.545 544.945 618.275 ;
      RECT 545.245 617.545 545.445 618.275 ;
      RECT 545.745 617.545 545.945 618.275 ;
      RECT 546.24 617.545 546.44 618.275 ;
      RECT 547.06 617.545 547.26 618.275 ;
      RECT 548.315 0.17 549.085 0.43 ;
      RECT 548.825 0.17 549.085 8.7 ;
      RECT 548.315 0.17 548.575 16.7 ;
      RECT 547.555 617.545 547.755 618.275 ;
      RECT 548.055 617.545 548.255 618.275 ;
      RECT 548.555 617.545 548.755 618.275 ;
      RECT 549.05 617.545 549.25 618.275 ;
      RECT 549.335 0.3 549.595 4.63 ;
      RECT 549.87 617.545 550.07 618.275 ;
      RECT 550.355 0.17 551.125 0.43 ;
      RECT 550.865 0.17 551.125 8.7 ;
      RECT 550.355 0.17 550.615 16.7 ;
      RECT 549.845 0.3 550.105 4.63 ;
      RECT 550.365 617.545 550.565 618.275 ;
      RECT 550.865 617.545 551.065 618.275 ;
      RECT 551.365 617.545 551.565 618.275 ;
      RECT 551.86 617.545 552.06 618.275 ;
      RECT 552.68 617.545 552.88 618.275 ;
      RECT 553.175 617.545 553.375 618.275 ;
      RECT 553.675 617.545 553.875 618.275 ;
      RECT 554.175 617.545 554.375 618.275 ;
      RECT 554.67 617.545 554.87 618.275 ;
      RECT 555.49 617.545 555.69 618.275 ;
      RECT 555.985 617.545 556.185 618.275 ;
      RECT 556.485 617.545 556.685 618.275 ;
      RECT 556.985 617.545 557.185 618.275 ;
      RECT 557.085 0.3 557.345 4.63 ;
      RECT 558.105 0.165 558.875 0.425 ;
      RECT 558.105 0.165 558.365 8.825 ;
      RECT 558.615 0.165 558.875 8.825 ;
      RECT 557.48 617.545 557.68 618.275 ;
      RECT 557.595 0.3 557.855 4.63 ;
      RECT 558.3 617.545 558.5 618.275 ;
      RECT 558.795 617.545 558.995 618.275 ;
      RECT 559.295 617.545 559.495 618.275 ;
      RECT 559.535 0.52 559.795 4.5 ;
      RECT 559.795 617.545 559.995 618.275 ;
      RECT 560.29 617.545 560.49 618.275 ;
      RECT 561.11 617.545 561.31 618.275 ;
      RECT 561.605 617.545 561.805 618.275 ;
      RECT 562.105 617.545 562.305 618.275 ;
      RECT 562.605 617.545 562.805 618.275 ;
      RECT 563.1 617.545 563.3 618.275 ;
      RECT 563.92 617.545 564.12 618.275 ;
      RECT 564.415 617.545 564.615 618.275 ;
      RECT 564.915 617.545 565.115 618.275 ;
      RECT 565.415 617.545 565.615 618.275 ;
      RECT 565.91 617.545 566.11 618.275 ;
      RECT 566.73 617.545 566.93 618.275 ;
      RECT 567.225 617.545 567.425 618.275 ;
      RECT 567.725 617.545 567.925 618.275 ;
      RECT 568.225 617.545 568.425 618.275 ;
      RECT 568.72 617.545 568.92 618.275 ;
      RECT 569.54 617.545 569.74 618.275 ;
      RECT 570.035 617.545 570.235 618.275 ;
      RECT 570.535 617.545 570.735 618.275 ;
      RECT 571.035 617.545 571.235 618.275 ;
      RECT 571.53 617.545 571.73 618.275 ;
      RECT 572.35 617.545 572.55 618.275 ;
      RECT 573.305 0.16 574.075 0.42 ;
      RECT 573.815 0.16 574.075 4.63 ;
      RECT 573.305 0.16 573.565 8.82 ;
      RECT 572.845 617.545 573.045 618.275 ;
      RECT 573.345 617.545 573.545 618.275 ;
      RECT 573.845 617.545 574.045 618.275 ;
      RECT 574.34 617.545 574.54 618.275 ;
      RECT 574.325 0.3 574.585 4.63 ;
      RECT 574.835 0.3 575.095 4.63 ;
      RECT 575.16 617.545 575.36 618.275 ;
      RECT 575.655 617.545 575.855 618.275 ;
      RECT 576.155 617.545 576.355 618.275 ;
      RECT 577.84 0.16 578.61 0.42 ;
      RECT 577.84 0.16 578.1 8.82 ;
      RECT 578.35 0.16 578.61 8.82 ;
      RECT 576.655 617.545 576.855 618.275 ;
      RECT 577.15 617.545 577.35 618.275 ;
      RECT 577.97 617.545 578.17 618.275 ;
      RECT 578.465 617.545 578.665 618.275 ;
      RECT 578.86 0.3 579.12 4.63 ;
      RECT 578.965 617.545 579.165 618.275 ;
      RECT 579.37 0.3 579.63 4.63 ;
      RECT 579.465 617.545 579.665 618.275 ;
      RECT 579.96 617.545 580.16 618.275 ;
      RECT 580.375 0.52 580.635 10.655 ;
      RECT 580.78 617.545 580.98 618.275 ;
      RECT 581.275 617.545 581.475 618.275 ;
      RECT 581.31 0.52 581.57 4.5 ;
      RECT 581.775 617.545 581.975 618.275 ;
      RECT 582.275 617.545 582.475 618.275 ;
      RECT 582.77 617.545 582.97 618.275 ;
      RECT 584.015 0.165 584.785 0.425 ;
      RECT 584.015 0.165 584.275 8.825 ;
      RECT 584.525 0.165 584.785 8.825 ;
      RECT 583.59 617.545 583.79 618.275 ;
      RECT 584.085 617.545 584.285 618.275 ;
      RECT 584.585 617.545 584.785 618.275 ;
      RECT 585.085 617.545 585.285 618.275 ;
      RECT 585.035 0.3 585.295 4.63 ;
      RECT 585.58 617.545 585.78 618.275 ;
      RECT 585.545 0.3 585.805 8.23 ;
      RECT 586.4 617.545 586.6 618.275 ;
      RECT 586.895 617.545 587.095 618.275 ;
      RECT 587.31 0.52 587.57 7.94 ;
      RECT 587.395 617.545 587.595 618.275 ;
      RECT 587.895 617.545 588.095 618.275 ;
      RECT 588.39 617.545 588.59 618.275 ;
      RECT 588.84 0.52 589.1 10.655 ;
      RECT 589.705 0.17 590.475 0.43 ;
      RECT 590.215 0.17 590.475 11.38 ;
      RECT 589.705 0.17 589.965 16.7 ;
      RECT 589.21 617.545 589.41 618.275 ;
      RECT 589.705 617.545 589.905 618.275 ;
      RECT 590.205 617.545 590.405 618.275 ;
      RECT 590.705 617.545 590.905 618.275 ;
      RECT 591.2 617.545 591.4 618.275 ;
      RECT 592.02 617.545 592.22 618.275 ;
      RECT 593.275 0.17 594.045 0.43 ;
      RECT 593.785 0.17 594.045 8.7 ;
      RECT 593.275 0.17 593.535 16.7 ;
      RECT 592.515 617.545 592.715 618.275 ;
      RECT 593.015 617.545 593.215 618.275 ;
      RECT 593.515 617.545 593.715 618.275 ;
      RECT 594.01 617.545 594.21 618.275 ;
      RECT 594.295 0.3 594.555 4.63 ;
      RECT 594.83 617.545 595.03 618.275 ;
      RECT 595.315 0.17 596.085 0.43 ;
      RECT 595.825 0.17 596.085 8.7 ;
      RECT 595.315 0.17 595.575 16.7 ;
      RECT 594.805 0.3 595.065 4.63 ;
      RECT 595.325 617.545 595.525 618.275 ;
      RECT 595.825 617.545 596.025 618.275 ;
      RECT 596.325 617.545 596.525 618.275 ;
      RECT 596.82 617.545 597.02 618.275 ;
      RECT 597.64 617.545 597.84 618.275 ;
      RECT 598.135 617.545 598.335 618.275 ;
      RECT 598.635 617.545 598.835 618.275 ;
      RECT 599.135 617.545 599.335 618.275 ;
      RECT 599.63 617.545 599.83 618.275 ;
      RECT 600.45 617.545 600.65 618.275 ;
      RECT 600.945 617.545 601.145 618.275 ;
      RECT 601.445 617.545 601.645 618.275 ;
      RECT 601.945 617.545 602.145 618.275 ;
      RECT 602.045 0.3 602.305 4.63 ;
      RECT 603.065 0.165 603.835 0.425 ;
      RECT 603.065 0.165 603.325 8.825 ;
      RECT 603.575 0.165 603.835 8.825 ;
      RECT 602.44 617.545 602.64 618.275 ;
      RECT 602.555 0.3 602.815 4.63 ;
      RECT 603.26 617.545 603.46 618.275 ;
      RECT 603.755 617.545 603.955 618.275 ;
      RECT 604.255 617.545 604.455 618.275 ;
      RECT 604.495 0.52 604.755 4.5 ;
      RECT 604.755 617.545 604.955 618.275 ;
      RECT 605.25 617.545 605.45 618.275 ;
      RECT 606.07 617.545 606.27 618.275 ;
      RECT 606.565 617.545 606.765 618.275 ;
      RECT 607.065 617.545 607.265 618.275 ;
      RECT 607.565 617.545 607.765 618.275 ;
      RECT 608.06 617.545 608.26 618.275 ;
      RECT 608.88 617.545 609.08 618.275 ;
      RECT 609.375 617.545 609.575 618.275 ;
      RECT 609.875 617.545 610.075 618.275 ;
      RECT 610.375 617.545 610.575 618.275 ;
      RECT 610.87 617.545 611.07 618.275 ;
      RECT 611.69 617.545 611.89 618.275 ;
      RECT 612.185 617.545 612.385 618.275 ;
      RECT 612.685 617.545 612.885 618.275 ;
      RECT 613.185 617.545 613.385 618.275 ;
      RECT 613.68 617.545 613.88 618.275 ;
      RECT 614.5 617.545 614.7 618.275 ;
      RECT 614.995 617.545 615.195 618.275 ;
      RECT 615.495 617.545 615.695 618.275 ;
      RECT 615.995 617.545 616.195 618.275 ;
      RECT 616.49 617.545 616.69 618.275 ;
      RECT 617.31 617.545 617.51 618.275 ;
      RECT 618.265 0.16 619.035 0.42 ;
      RECT 618.775 0.16 619.035 4.63 ;
      RECT 618.265 0.16 618.525 8.82 ;
      RECT 617.805 617.545 618.005 618.275 ;
      RECT 618.305 617.545 618.505 618.275 ;
      RECT 618.805 617.545 619.005 618.275 ;
      RECT 619.3 617.545 619.5 618.275 ;
      RECT 619.285 0.3 619.545 4.63 ;
      RECT 619.795 0.3 620.055 4.63 ;
      RECT 620.12 617.545 620.32 618.275 ;
      RECT 620.615 617.545 620.815 618.275 ;
      RECT 621.115 617.545 621.315 618.275 ;
      RECT 622.8 0.16 623.57 0.42 ;
      RECT 622.8 0.16 623.06 8.82 ;
      RECT 623.31 0.16 623.57 8.82 ;
      RECT 621.615 617.545 621.815 618.275 ;
      RECT 622.11 617.545 622.31 618.275 ;
      RECT 622.93 617.545 623.13 618.275 ;
      RECT 623.425 617.545 623.625 618.275 ;
      RECT 623.82 0.3 624.08 4.63 ;
      RECT 623.925 617.545 624.125 618.275 ;
      RECT 624.33 0.3 624.59 4.63 ;
      RECT 624.425 617.545 624.625 618.275 ;
      RECT 624.92 617.545 625.12 618.275 ;
      RECT 625.335 0.52 625.595 10.655 ;
      RECT 625.74 617.545 625.94 618.275 ;
      RECT 626.235 617.545 626.435 618.275 ;
      RECT 626.27 0.52 626.53 4.5 ;
      RECT 626.735 617.545 626.935 618.275 ;
      RECT 627.235 617.545 627.435 618.275 ;
      RECT 627.73 617.545 627.93 618.275 ;
      RECT 628.975 0.165 629.745 0.425 ;
      RECT 628.975 0.165 629.235 8.825 ;
      RECT 629.485 0.165 629.745 8.825 ;
      RECT 628.55 617.545 628.75 618.275 ;
      RECT 629.045 617.545 629.245 618.275 ;
      RECT 629.545 617.545 629.745 618.275 ;
      RECT 630.045 617.545 630.245 618.275 ;
      RECT 629.995 0.3 630.255 4.63 ;
      RECT 630.54 617.545 630.74 618.275 ;
      RECT 630.505 0.3 630.765 8.23 ;
      RECT 631.36 617.545 631.56 618.275 ;
      RECT 631.855 617.545 632.055 618.275 ;
      RECT 632.27 0.52 632.53 7.94 ;
      RECT 632.355 617.545 632.555 618.275 ;
      RECT 632.855 617.545 633.055 618.275 ;
      RECT 633.35 617.545 633.55 618.275 ;
      RECT 633.8 0.52 634.06 10.655 ;
      RECT 634.665 0.17 635.435 0.43 ;
      RECT 635.175 0.17 635.435 11.38 ;
      RECT 634.665 0.17 634.925 16.7 ;
      RECT 634.17 617.545 634.37 618.275 ;
      RECT 634.665 617.545 634.865 618.275 ;
      RECT 635.165 617.545 635.365 618.275 ;
      RECT 635.665 617.545 635.865 618.275 ;
      RECT 636.16 617.545 636.36 618.275 ;
      RECT 636.98 617.545 637.18 618.275 ;
      RECT 638.235 0.17 639.005 0.43 ;
      RECT 638.745 0.17 639.005 8.7 ;
      RECT 638.235 0.17 638.495 16.7 ;
      RECT 637.475 617.545 637.675 618.275 ;
      RECT 637.975 617.545 638.175 618.275 ;
      RECT 638.475 617.545 638.675 618.275 ;
      RECT 638.97 617.545 639.17 618.275 ;
      RECT 639.255 0.3 639.515 4.63 ;
      RECT 639.79 617.545 639.99 618.275 ;
      RECT 640.275 0.17 641.045 0.43 ;
      RECT 640.785 0.17 641.045 8.7 ;
      RECT 640.275 0.17 640.535 16.7 ;
      RECT 639.765 0.3 640.025 4.63 ;
      RECT 640.285 617.545 640.485 618.275 ;
      RECT 640.785 617.545 640.985 618.275 ;
      RECT 641.285 617.545 641.485 618.275 ;
      RECT 641.78 617.545 641.98 618.275 ;
      RECT 642.6 617.545 642.8 618.275 ;
      RECT 643.095 617.545 643.295 618.275 ;
      RECT 643.595 617.545 643.795 618.275 ;
      RECT 644.095 617.545 644.295 618.275 ;
      RECT 644.59 617.545 644.79 618.275 ;
      RECT 645.41 617.545 645.61 618.275 ;
      RECT 645.905 617.545 646.105 618.275 ;
      RECT 646.405 617.545 646.605 618.275 ;
      RECT 646.905 617.545 647.105 618.275 ;
      RECT 647.005 0.3 647.265 4.63 ;
      RECT 648.025 0.165 648.795 0.425 ;
      RECT 648.025 0.165 648.285 8.825 ;
      RECT 648.535 0.165 648.795 8.825 ;
      RECT 647.4 617.545 647.6 618.275 ;
      RECT 647.515 0.3 647.775 4.63 ;
      RECT 648.22 617.545 648.42 618.275 ;
      RECT 648.715 617.545 648.915 618.275 ;
      RECT 649.215 617.545 649.415 618.275 ;
      RECT 649.455 0.52 649.715 4.5 ;
      RECT 649.715 617.545 649.915 618.275 ;
      RECT 650.21 617.545 650.41 618.275 ;
      RECT 651.03 617.545 651.23 618.275 ;
      RECT 651.525 617.545 651.725 618.275 ;
      RECT 652.025 617.545 652.225 618.275 ;
      RECT 652.525 617.545 652.725 618.275 ;
      RECT 653.02 617.545 653.22 618.275 ;
      RECT 653.84 617.545 654.04 618.275 ;
      RECT 654.335 617.545 654.535 618.275 ;
      RECT 654.835 617.545 655.035 618.275 ;
      RECT 655.335 617.545 655.535 618.275 ;
      RECT 655.83 617.545 656.03 618.275 ;
      RECT 656.65 617.545 656.85 618.275 ;
      RECT 657.145 617.545 657.345 618.275 ;
      RECT 657.645 617.545 657.845 618.275 ;
      RECT 658.145 617.545 658.345 618.275 ;
      RECT 658.64 617.545 658.84 618.275 ;
      RECT 659.46 617.545 659.66 618.275 ;
      RECT 659.955 617.545 660.155 618.275 ;
      RECT 660.455 617.545 660.655 618.275 ;
      RECT 660.955 617.545 661.155 618.275 ;
      RECT 661.45 617.545 661.65 618.275 ;
      RECT 662.27 617.545 662.47 618.275 ;
      RECT 663.225 0.16 663.995 0.42 ;
      RECT 663.735 0.16 663.995 4.63 ;
      RECT 663.225 0.16 663.485 8.82 ;
      RECT 662.765 617.545 662.965 618.275 ;
      RECT 663.265 617.545 663.465 618.275 ;
      RECT 663.765 617.545 663.965 618.275 ;
      RECT 664.26 617.545 664.46 618.275 ;
      RECT 664.245 0.3 664.505 4.63 ;
      RECT 664.755 0.3 665.015 4.63 ;
      RECT 665.08 617.545 665.28 618.275 ;
      RECT 665.575 617.545 665.775 618.275 ;
      RECT 666.075 617.545 666.275 618.275 ;
      RECT 667.76 0.16 668.53 0.42 ;
      RECT 667.76 0.16 668.02 8.82 ;
      RECT 668.27 0.16 668.53 8.82 ;
      RECT 666.575 617.545 666.775 618.275 ;
      RECT 667.07 617.545 667.27 618.275 ;
      RECT 667.89 617.545 668.09 618.275 ;
      RECT 668.385 617.545 668.585 618.275 ;
      RECT 668.78 0.3 669.04 4.63 ;
      RECT 668.885 617.545 669.085 618.275 ;
      RECT 669.29 0.3 669.55 4.63 ;
      RECT 669.385 617.545 669.585 618.275 ;
      RECT 669.88 617.545 670.08 618.275 ;
      RECT 670.295 0.52 670.555 10.655 ;
      RECT 670.7 617.545 670.9 618.275 ;
      RECT 671.195 617.545 671.395 618.275 ;
      RECT 671.23 0.52 671.49 4.5 ;
      RECT 671.695 617.545 671.895 618.275 ;
      RECT 672.195 617.545 672.395 618.275 ;
      RECT 672.69 617.545 672.89 618.275 ;
      RECT 673.935 0.165 674.705 0.425 ;
      RECT 673.935 0.165 674.195 8.825 ;
      RECT 674.445 0.165 674.705 8.825 ;
      RECT 673.51 617.545 673.71 618.275 ;
      RECT 674.005 617.545 674.205 618.275 ;
      RECT 674.505 617.545 674.705 618.275 ;
      RECT 675.005 617.545 675.205 618.275 ;
      RECT 674.955 0.3 675.215 4.63 ;
      RECT 675.5 617.545 675.7 618.275 ;
      RECT 675.465 0.3 675.725 8.23 ;
      RECT 676.32 617.545 676.52 618.275 ;
      RECT 676.815 617.545 677.015 618.275 ;
      RECT 677.23 0.52 677.49 7.94 ;
      RECT 677.315 617.545 677.515 618.275 ;
      RECT 677.815 617.545 678.015 618.275 ;
      RECT 678.31 617.545 678.51 618.275 ;
      RECT 678.76 0.52 679.02 10.655 ;
      RECT 679.625 0.17 680.395 0.43 ;
      RECT 680.135 0.17 680.395 11.38 ;
      RECT 679.625 0.17 679.885 16.7 ;
      RECT 679.13 617.545 679.33 618.275 ;
      RECT 679.625 617.545 679.825 618.275 ;
      RECT 680.125 617.545 680.325 618.275 ;
      RECT 680.625 617.545 680.825 618.275 ;
      RECT 681.12 617.545 681.32 618.275 ;
      RECT 681.94 617.545 682.14 618.275 ;
      RECT 683.195 0.17 683.965 0.43 ;
      RECT 683.705 0.17 683.965 8.7 ;
      RECT 683.195 0.17 683.455 16.7 ;
      RECT 682.435 617.545 682.635 618.275 ;
      RECT 682.935 617.545 683.135 618.275 ;
      RECT 683.435 617.545 683.635 618.275 ;
      RECT 683.93 617.545 684.13 618.275 ;
      RECT 684.215 0.3 684.475 4.63 ;
      RECT 684.75 617.545 684.95 618.275 ;
      RECT 685.235 0.17 686.005 0.43 ;
      RECT 685.745 0.17 686.005 8.7 ;
      RECT 685.235 0.17 685.495 16.7 ;
      RECT 684.725 0.3 684.985 4.63 ;
      RECT 685.245 617.545 685.445 618.275 ;
      RECT 685.745 617.545 685.945 618.275 ;
      RECT 686.245 617.545 686.445 618.275 ;
      RECT 686.74 617.545 686.94 618.275 ;
      RECT 687.56 617.545 687.76 618.275 ;
      RECT 688.055 617.545 688.255 618.275 ;
      RECT 688.555 617.545 688.755 618.275 ;
      RECT 689.055 617.545 689.255 618.275 ;
      RECT 689.55 617.545 689.75 618.275 ;
      RECT 690.37 617.545 690.57 618.275 ;
      RECT 690.865 617.545 691.065 618.275 ;
      RECT 691.365 617.545 691.565 618.275 ;
      RECT 691.865 617.545 692.065 618.275 ;
      RECT 691.965 0.3 692.225 4.63 ;
      RECT 692.985 0.165 693.755 0.425 ;
      RECT 692.985 0.165 693.245 8.825 ;
      RECT 693.495 0.165 693.755 8.825 ;
      RECT 692.36 617.545 692.56 618.275 ;
      RECT 692.475 0.3 692.735 4.63 ;
      RECT 693.18 617.545 693.38 618.275 ;
      RECT 693.675 617.545 693.875 618.275 ;
      RECT 694.175 617.545 694.375 618.275 ;
      RECT 694.415 0.52 694.675 4.5 ;
      RECT 694.675 617.545 694.875 618.275 ;
      RECT 695.17 617.545 695.37 618.275 ;
      RECT 695.99 617.545 696.19 618.275 ;
      RECT 696.485 617.545 696.685 618.275 ;
      RECT 696.985 617.545 697.185 618.275 ;
      RECT 697.485 617.545 697.685 618.275 ;
      RECT 697.98 617.545 698.18 618.275 ;
      RECT 698.8 617.545 699 618.275 ;
      RECT 699.295 617.545 699.495 618.275 ;
      RECT 699.795 617.545 699.995 618.275 ;
      RECT 700.295 617.545 700.495 618.275 ;
      RECT 700.79 617.545 700.99 618.275 ;
      RECT 701.61 617.545 701.81 618.275 ;
      RECT 702.105 617.545 702.305 618.275 ;
      RECT 702.605 617.545 702.805 618.275 ;
      RECT 703.105 617.545 703.305 618.275 ;
      RECT 703.6 617.545 703.8 618.275 ;
      RECT 704.42 617.545 704.62 618.275 ;
      RECT 704.915 617.545 705.115 618.275 ;
      RECT 705.415 617.545 705.615 618.275 ;
      RECT 705.915 617.545 706.115 618.275 ;
      RECT 706.41 617.545 706.61 618.275 ;
      RECT 707.23 617.545 707.43 618.275 ;
      RECT 708.185 0.16 708.955 0.42 ;
      RECT 708.695 0.16 708.955 4.63 ;
      RECT 708.185 0.16 708.445 8.82 ;
      RECT 707.725 617.545 707.925 618.275 ;
      RECT 708.225 617.545 708.425 618.275 ;
      RECT 708.725 617.545 708.925 618.275 ;
      RECT 709.22 617.545 709.42 618.275 ;
      RECT 709.205 0.3 709.465 4.63 ;
      RECT 709.715 0.3 709.975 4.63 ;
      RECT 710.04 617.545 710.24 618.275 ;
      RECT 710.535 617.545 710.735 618.275 ;
      RECT 711.035 617.545 711.235 618.275 ;
      RECT 712.72 0.16 713.49 0.42 ;
      RECT 712.72 0.16 712.98 8.82 ;
      RECT 713.23 0.16 713.49 8.82 ;
      RECT 711.535 617.545 711.735 618.275 ;
      RECT 712.03 617.545 712.23 618.275 ;
      RECT 712.85 617.545 713.05 618.275 ;
      RECT 713.345 617.545 713.545 618.275 ;
      RECT 713.74 0.3 714 4.63 ;
      RECT 713.845 617.545 714.045 618.275 ;
      RECT 714.25 0.3 714.51 4.63 ;
      RECT 714.345 617.545 714.545 618.275 ;
      RECT 714.84 617.545 715.04 618.275 ;
      RECT 715.255 0.52 715.515 10.655 ;
      RECT 715.66 617.545 715.86 618.275 ;
      RECT 716.155 617.545 716.355 618.275 ;
      RECT 716.19 0.52 716.45 4.5 ;
      RECT 716.655 617.545 716.855 618.275 ;
      RECT 717.155 617.545 717.355 618.275 ;
      RECT 717.65 617.545 717.85 618.275 ;
      RECT 718.895 0.165 719.665 0.425 ;
      RECT 718.895 0.165 719.155 8.825 ;
      RECT 719.405 0.165 719.665 8.825 ;
      RECT 718.47 617.545 718.67 618.275 ;
      RECT 718.965 617.545 719.165 618.275 ;
      RECT 719.465 617.545 719.665 618.275 ;
      RECT 719.965 617.545 720.165 618.275 ;
      RECT 719.915 0.3 720.175 4.63 ;
      RECT 720.46 617.545 720.66 618.275 ;
      RECT 720.425 0.3 720.685 8.23 ;
      RECT 721.28 617.545 721.48 618.275 ;
      RECT 723.995 0.17 724.765 0.43 ;
      RECT 723.995 0.17 724.255 34.45 ;
      RECT 724.505 0.17 724.765 34.45 ;
      RECT 722.275 617.545 722.475 618.275 ;
      RECT 722.975 0.3 723.235 35.29 ;
      RECT 723.485 0.3 723.745 35.29 ;
      RECT 725.015 0.3 725.275 35.29 ;
      RECT 725.525 0.3 725.785 35.29 ;
      RECT 730.115 0.17 730.885 0.43 ;
      RECT 730.115 0.17 730.375 34.03 ;
      RECT 730.625 0.17 730.885 34.03 ;
      RECT 726.035 0.3 726.295 34.03 ;
      RECT 729.095 0.3 729.355 35.29 ;
      RECT 729.605 0.3 729.865 35.29 ;
      RECT 731.135 0.3 731.395 35.29 ;
      RECT 734.195 0.17 734.965 0.43 ;
      RECT 734.195 0.17 734.455 36.945 ;
      RECT 734.705 0.17 734.965 36.945 ;
      RECT 731.645 0.3 731.905 35.29 ;
      RECT 732.155 0.3 732.415 34.03 ;
      RECT 736.235 0.17 737.005 0.43 ;
      RECT 736.235 0.17 736.495 36.945 ;
      RECT 736.745 0.17 737.005 36.945 ;
      RECT 732.665 0.3 732.925 2.225 ;
      RECT 735.215 0.3 735.475 37.365 ;
      RECT 738.275 0.17 739.045 0.43 ;
      RECT 738.275 0.17 738.535 36.945 ;
      RECT 738.785 0.17 739.045 36.945 ;
      RECT 735.725 0.3 735.985 37.365 ;
      RECT 737.255 0.3 737.515 37.365 ;
      RECT 740.98 0 741.24 4.94 ;
      RECT 740.98 4.68 741.75 4.94 ;
      RECT 741.49 4.68 741.75 12.9 ;
      RECT 741.49 0.52 741.75 1.78 ;
      RECT 741.49 1.52 742.26 1.78 ;
      RECT 742 1.52 742.26 12.9 ;
      RECT 737.765 0.3 738.025 37.365 ;
      RECT 742 0.59 742.77 1.27 ;
      RECT 742.51 0.59 742.77 7.965 ;
      RECT 739.295 0.3 739.555 37.365 ;
      RECT 739.805 0.3 740.065 37.365 ;
      RECT 743.02 0.52 743.28 12.9 ;
      RECT 743.53 0 743.79 12.9 ;
      RECT 744.04 0.52 744.3 12.9 ;
      RECT 744.55 0.52 744.81 12.9 ;
      RECT 745.06 0.52 745.32 12.9 ;
      RECT 745.57 0.52 745.83 12.9 ;
      RECT 747.1 0.59 747.87 1.27 ;
      RECT 748.12 0.17 748.89 0.43 ;
      RECT 748.12 0.17 748.38 2.085 ;
      RECT 748.63 0.17 748.89 9 ;
      RECT 747.1 0.59 747.36 7.545 ;
      RECT 746.08 0.52 746.34 8.565 ;
      RECT 746.59 0.52 746.85 8.055 ;
      RECT 752.71 0.52 752.97 6.59 ;
      RECT 754.24 0.52 754.5 6.305 ;
      RECT 754.24 6.045 755.21 6.305 ;
      RECT 753.22 0.52 753.48 2.23 ;
      RECT 754.75 0.52 755.01 2.955 ;
      RECT 755.77 0.52 756.03 12.9 ;
      RECT 756.28 0.52 756.54 12.9 ;
      RECT 757.81 0.52 758.07 6.29 ;
      RECT 757.3 6.045 758.07 6.29 ;
      RECT 756.79 0.52 757.05 6.745 ;
      RECT 759.34 0.52 759.6 6.59 ;
      RECT 758.695 6.33 759.6 6.59 ;
      RECT 757.3 0.52 757.56 2.955 ;
      RECT 758.83 0.52 759.09 2.67 ;
      RECT 760.36 0.52 760.62 12.9 ;
      RECT 760.87 0.52 761.13 12.9 ;
      RECT 762.4 0.575 762.66 7.965 ;
      RECT 762.91 0.52 763.17 12.9 ;
      RECT 763.42 0.52 763.68 12.9 ;
      RECT 763.93 0.52 764.19 12.9 ;
      RECT 764.44 0.52 764.7 12.9 ;
      RECT 764.95 0.52 765.21 12.9 ;
      RECT 765.46 0.52 765.72 12.9 ;
      RECT 765.97 0.52 766.23 12.9 ;
      RECT 766.48 0.52 766.74 12.9 ;
      RECT 768.01 0.59 768.78 1.27 ;
      RECT 768.01 0.59 768.27 8.83 ;
      RECT 766.99 0.52 767.25 12.9 ;
      RECT 767.5 0.52 767.76 12.9 ;
      RECT 769.03 0.52 769.29 12.9 ;
      RECT 769.54 0.52 769.8 12.9 ;
      RECT 776.68 0.17 777.45 0.43 ;
      RECT 776.68 0.17 776.94 13.845 ;
      RECT 777.19 0.17 777.45 13.845 ;
      RECT 778.72 0.17 779.49 0.43 ;
      RECT 778.72 0.17 778.98 2.11 ;
      RECT 779.23 0.17 779.49 2.11 ;
      RECT 774.13 0.52 774.39 3.61 ;
      RECT 774.64 0.52 774.9 4.12 ;
      RECT 781.115 0.17 781.885 0.43 ;
      RECT 781.115 0.17 781.375 36.945 ;
      RECT 781.625 0.17 781.885 36.945 ;
      RECT 776.17 0.52 776.43 15.16 ;
      RECT 780.095 0.3 780.355 37.365 ;
      RECT 783.155 0.17 783.925 0.43 ;
      RECT 783.155 0.17 783.415 36.945 ;
      RECT 783.665 0.17 783.925 36.945 ;
      RECT 780.605 0.3 780.865 37.365 ;
      RECT 782.135 0.3 782.395 37.365 ;
      RECT 785.195 0.17 785.965 0.43 ;
      RECT 785.195 0.17 785.455 36.945 ;
      RECT 785.705 0.17 785.965 36.945 ;
      RECT 782.645 0.3 782.905 37.365 ;
      RECT 784.175 0.3 784.435 37.365 ;
      RECT 784.685 0.3 784.945 37.365 ;
      RECT 787.235 0.3 787.495 2.225 ;
      RECT 789.275 0.17 790.045 0.43 ;
      RECT 789.275 0.17 789.535 34.03 ;
      RECT 789.785 0.17 790.045 34.03 ;
      RECT 787.745 0.3 788.005 34.03 ;
      RECT 788.255 0.3 788.515 35.29 ;
      RECT 788.765 0.3 789.025 35.29 ;
      RECT 790.295 0.3 790.555 35.29 ;
      RECT 790.805 0.3 791.065 35.29 ;
      RECT 795.395 0.17 796.165 0.43 ;
      RECT 795.395 0.17 795.655 34.45 ;
      RECT 795.905 0.17 796.165 34.45 ;
      RECT 793.865 0.3 794.125 34.03 ;
      RECT 794.375 0.3 794.635 35.29 ;
      RECT 794.885 0.3 795.145 35.29 ;
      RECT 796.415 0.3 796.675 35.29 ;
      RECT 796.925 0.3 797.185 35.29 ;
      RECT 797.685 617.545 797.885 618.275 ;
      RECT 798.68 617.545 798.88 618.275 ;
      RECT 799.5 617.545 799.7 618.275 ;
      RECT 799.475 0.3 799.735 8.23 ;
      RECT 799.995 617.545 800.195 618.275 ;
      RECT 800.495 0.165 801.265 0.425 ;
      RECT 800.495 0.165 800.755 8.825 ;
      RECT 801.005 0.165 801.265 8.825 ;
      RECT 799.985 0.3 800.245 4.63 ;
      RECT 800.495 617.545 800.695 618.275 ;
      RECT 800.995 617.545 801.195 618.275 ;
      RECT 801.49 617.545 801.69 618.275 ;
      RECT 802.31 617.545 802.51 618.275 ;
      RECT 802.805 617.545 803.005 618.275 ;
      RECT 803.305 617.545 803.505 618.275 ;
      RECT 803.71 0.52 803.97 4.5 ;
      RECT 803.805 617.545 804.005 618.275 ;
      RECT 804.3 617.545 804.5 618.275 ;
      RECT 804.645 0.52 804.905 10.655 ;
      RECT 805.12 617.545 805.32 618.275 ;
      RECT 805.615 617.545 805.815 618.275 ;
      RECT 805.65 0.3 805.91 4.63 ;
      RECT 806.115 617.545 806.315 618.275 ;
      RECT 806.67 0.16 807.44 0.42 ;
      RECT 806.67 0.16 806.93 8.82 ;
      RECT 807.18 0.16 807.44 8.82 ;
      RECT 806.16 0.3 806.42 4.63 ;
      RECT 806.615 617.545 806.815 618.275 ;
      RECT 807.11 617.545 807.31 618.275 ;
      RECT 807.93 617.545 808.13 618.275 ;
      RECT 808.425 617.545 808.625 618.275 ;
      RECT 808.925 617.545 809.125 618.275 ;
      RECT 809.425 617.545 809.625 618.275 ;
      RECT 809.92 617.545 810.12 618.275 ;
      RECT 810.185 0.3 810.445 4.63 ;
      RECT 810.74 617.545 810.94 618.275 ;
      RECT 811.205 0.16 811.975 0.42 ;
      RECT 811.205 0.16 811.465 4.63 ;
      RECT 811.715 0.16 811.975 8.82 ;
      RECT 810.695 0.3 810.955 4.63 ;
      RECT 811.235 617.545 811.435 618.275 ;
      RECT 811.735 617.545 811.935 618.275 ;
      RECT 812.235 617.545 812.435 618.275 ;
      RECT 812.73 617.545 812.93 618.275 ;
      RECT 813.55 617.545 813.75 618.275 ;
      RECT 814.045 617.545 814.245 618.275 ;
      RECT 814.545 617.545 814.745 618.275 ;
      RECT 815.045 617.545 815.245 618.275 ;
      RECT 815.54 617.545 815.74 618.275 ;
      RECT 816.36 617.545 816.56 618.275 ;
      RECT 816.855 617.545 817.055 618.275 ;
      RECT 817.355 617.545 817.555 618.275 ;
      RECT 817.855 617.545 818.055 618.275 ;
      RECT 818.35 617.545 818.55 618.275 ;
      RECT 819.17 617.545 819.37 618.275 ;
      RECT 819.665 617.545 819.865 618.275 ;
      RECT 820.165 617.545 820.365 618.275 ;
      RECT 820.665 617.545 820.865 618.275 ;
      RECT 821.16 617.545 821.36 618.275 ;
      RECT 821.98 617.545 822.18 618.275 ;
      RECT 822.475 617.545 822.675 618.275 ;
      RECT 822.975 617.545 823.175 618.275 ;
      RECT 823.475 617.545 823.675 618.275 ;
      RECT 823.97 617.545 824.17 618.275 ;
      RECT 824.79 617.545 824.99 618.275 ;
      RECT 825.285 617.545 825.485 618.275 ;
      RECT 825.485 0.52 825.745 4.5 ;
      RECT 826.405 0.165 827.175 0.425 ;
      RECT 826.405 0.165 826.665 8.825 ;
      RECT 826.915 0.165 827.175 8.825 ;
      RECT 825.785 617.545 825.985 618.275 ;
      RECT 826.285 617.545 826.485 618.275 ;
      RECT 826.78 617.545 826.98 618.275 ;
      RECT 827.425 0.3 827.685 4.63 ;
      RECT 827.6 617.545 827.8 618.275 ;
      RECT 827.935 0.3 828.195 4.63 ;
      RECT 828.095 617.545 828.295 618.275 ;
      RECT 828.595 617.545 828.795 618.275 ;
      RECT 829.095 617.545 829.295 618.275 ;
      RECT 829.59 617.545 829.79 618.275 ;
      RECT 830.41 617.545 830.61 618.275 ;
      RECT 830.905 617.545 831.105 618.275 ;
      RECT 831.405 617.545 831.605 618.275 ;
      RECT 831.905 617.545 832.105 618.275 ;
      RECT 832.4 617.545 832.6 618.275 ;
      RECT 833.22 617.545 833.42 618.275 ;
      RECT 834.155 0.17 834.925 0.43 ;
      RECT 834.155 0.17 834.415 8.7 ;
      RECT 834.665 0.17 834.925 16.7 ;
      RECT 833.715 617.545 833.915 618.275 ;
      RECT 834.215 617.545 834.415 618.275 ;
      RECT 834.715 617.545 834.915 618.275 ;
      RECT 835.21 617.545 835.41 618.275 ;
      RECT 835.175 0.3 835.435 4.63 ;
      RECT 836.195 0.17 836.965 0.43 ;
      RECT 836.195 0.17 836.455 8.7 ;
      RECT 836.705 0.17 836.965 16.7 ;
      RECT 835.685 0.3 835.945 4.63 ;
      RECT 836.03 617.545 836.23 618.275 ;
      RECT 836.525 617.545 836.725 618.275 ;
      RECT 837.025 617.545 837.225 618.275 ;
      RECT 837.525 617.545 837.725 618.275 ;
      RECT 838.02 617.545 838.22 618.275 ;
      RECT 838.84 617.545 839.04 618.275 ;
      RECT 839.765 0.17 840.535 0.43 ;
      RECT 839.765 0.17 840.025 11.38 ;
      RECT 840.275 0.17 840.535 16.7 ;
      RECT 839.335 617.545 839.535 618.275 ;
      RECT 839.835 617.545 840.035 618.275 ;
      RECT 840.335 617.545 840.535 618.275 ;
      RECT 840.83 617.545 841.03 618.275 ;
      RECT 841.14 0.52 841.4 10.655 ;
      RECT 841.65 617.545 841.85 618.275 ;
      RECT 842.145 617.545 842.345 618.275 ;
      RECT 842.645 617.545 842.845 618.275 ;
      RECT 842.67 0.52 842.93 7.94 ;
      RECT 843.145 617.545 843.345 618.275 ;
      RECT 843.64 617.545 843.84 618.275 ;
      RECT 844.46 617.545 844.66 618.275 ;
      RECT 844.435 0.3 844.695 8.23 ;
      RECT 844.955 617.545 845.155 618.275 ;
      RECT 845.455 0.165 846.225 0.425 ;
      RECT 845.455 0.165 845.715 8.825 ;
      RECT 845.965 0.165 846.225 8.825 ;
      RECT 844.945 0.3 845.205 4.63 ;
      RECT 845.455 617.545 845.655 618.275 ;
      RECT 845.955 617.545 846.155 618.275 ;
      RECT 846.45 617.545 846.65 618.275 ;
      RECT 847.27 617.545 847.47 618.275 ;
      RECT 847.765 617.545 847.965 618.275 ;
      RECT 848.265 617.545 848.465 618.275 ;
      RECT 848.67 0.52 848.93 4.5 ;
      RECT 848.765 617.545 848.965 618.275 ;
      RECT 849.26 617.545 849.46 618.275 ;
      RECT 849.605 0.52 849.865 10.655 ;
      RECT 850.08 617.545 850.28 618.275 ;
      RECT 850.575 617.545 850.775 618.275 ;
      RECT 850.61 0.3 850.87 4.63 ;
      RECT 851.075 617.545 851.275 618.275 ;
      RECT 851.63 0.16 852.4 0.42 ;
      RECT 851.63 0.16 851.89 8.82 ;
      RECT 852.14 0.16 852.4 8.82 ;
      RECT 851.12 0.3 851.38 4.63 ;
      RECT 851.575 617.545 851.775 618.275 ;
      RECT 852.07 617.545 852.27 618.275 ;
      RECT 852.89 617.545 853.09 618.275 ;
      RECT 853.385 617.545 853.585 618.275 ;
      RECT 853.885 617.545 854.085 618.275 ;
      RECT 854.385 617.545 854.585 618.275 ;
      RECT 854.88 617.545 855.08 618.275 ;
      RECT 855.145 0.3 855.405 4.63 ;
      RECT 855.7 617.545 855.9 618.275 ;
      RECT 856.165 0.16 856.935 0.42 ;
      RECT 856.165 0.16 856.425 4.63 ;
      RECT 856.675 0.16 856.935 8.82 ;
      RECT 855.655 0.3 855.915 4.63 ;
      RECT 856.195 617.545 856.395 618.275 ;
      RECT 856.695 617.545 856.895 618.275 ;
      RECT 857.195 617.545 857.395 618.275 ;
      RECT 857.69 617.545 857.89 618.275 ;
      RECT 858.51 617.545 858.71 618.275 ;
      RECT 859.005 617.545 859.205 618.275 ;
      RECT 859.505 617.545 859.705 618.275 ;
      RECT 860.005 617.545 860.205 618.275 ;
      RECT 860.5 617.545 860.7 618.275 ;
      RECT 861.32 617.545 861.52 618.275 ;
      RECT 861.815 617.545 862.015 618.275 ;
      RECT 862.315 617.545 862.515 618.275 ;
      RECT 862.815 617.545 863.015 618.275 ;
      RECT 863.31 617.545 863.51 618.275 ;
      RECT 864.13 617.545 864.33 618.275 ;
      RECT 864.625 617.545 864.825 618.275 ;
      RECT 865.125 617.545 865.325 618.275 ;
      RECT 865.625 617.545 865.825 618.275 ;
      RECT 866.12 617.545 866.32 618.275 ;
      RECT 866.94 617.545 867.14 618.275 ;
      RECT 867.435 617.545 867.635 618.275 ;
      RECT 867.935 617.545 868.135 618.275 ;
      RECT 868.435 617.545 868.635 618.275 ;
      RECT 868.93 617.545 869.13 618.275 ;
      RECT 869.75 617.545 869.95 618.275 ;
      RECT 870.245 617.545 870.445 618.275 ;
      RECT 870.445 0.52 870.705 4.5 ;
      RECT 871.365 0.165 872.135 0.425 ;
      RECT 871.365 0.165 871.625 8.825 ;
      RECT 871.875 0.165 872.135 8.825 ;
      RECT 870.745 617.545 870.945 618.275 ;
      RECT 871.245 617.545 871.445 618.275 ;
      RECT 871.74 617.545 871.94 618.275 ;
      RECT 872.385 0.3 872.645 4.63 ;
      RECT 872.56 617.545 872.76 618.275 ;
      RECT 872.895 0.3 873.155 4.63 ;
      RECT 873.055 617.545 873.255 618.275 ;
      RECT 873.555 617.545 873.755 618.275 ;
      RECT 874.055 617.545 874.255 618.275 ;
      RECT 874.55 617.545 874.75 618.275 ;
      RECT 875.37 617.545 875.57 618.275 ;
      RECT 875.865 617.545 876.065 618.275 ;
      RECT 876.365 617.545 876.565 618.275 ;
      RECT 876.865 617.545 877.065 618.275 ;
      RECT 877.36 617.545 877.56 618.275 ;
      RECT 878.18 617.545 878.38 618.275 ;
      RECT 879.115 0.17 879.885 0.43 ;
      RECT 879.115 0.17 879.375 8.7 ;
      RECT 879.625 0.17 879.885 16.7 ;
      RECT 878.675 617.545 878.875 618.275 ;
      RECT 879.175 617.545 879.375 618.275 ;
      RECT 879.675 617.545 879.875 618.275 ;
      RECT 880.17 617.545 880.37 618.275 ;
      RECT 880.135 0.3 880.395 4.63 ;
      RECT 881.155 0.17 881.925 0.43 ;
      RECT 881.155 0.17 881.415 8.7 ;
      RECT 881.665 0.17 881.925 16.7 ;
      RECT 880.645 0.3 880.905 4.63 ;
      RECT 880.99 617.545 881.19 618.275 ;
      RECT 881.485 617.545 881.685 618.275 ;
      RECT 881.985 617.545 882.185 618.275 ;
      RECT 882.485 617.545 882.685 618.275 ;
      RECT 882.98 617.545 883.18 618.275 ;
      RECT 883.8 617.545 884 618.275 ;
      RECT 884.725 0.17 885.495 0.43 ;
      RECT 884.725 0.17 884.985 11.38 ;
      RECT 885.235 0.17 885.495 16.7 ;
      RECT 884.295 617.545 884.495 618.275 ;
      RECT 884.795 617.545 884.995 618.275 ;
      RECT 885.295 617.545 885.495 618.275 ;
      RECT 885.79 617.545 885.99 618.275 ;
      RECT 886.1 0.52 886.36 10.655 ;
      RECT 886.61 617.545 886.81 618.275 ;
      RECT 887.105 617.545 887.305 618.275 ;
      RECT 887.605 617.545 887.805 618.275 ;
      RECT 887.63 0.52 887.89 7.94 ;
      RECT 888.105 617.545 888.305 618.275 ;
      RECT 888.6 617.545 888.8 618.275 ;
      RECT 889.42 617.545 889.62 618.275 ;
      RECT 889.395 0.3 889.655 8.23 ;
      RECT 889.915 617.545 890.115 618.275 ;
      RECT 890.415 0.165 891.185 0.425 ;
      RECT 890.415 0.165 890.675 8.825 ;
      RECT 890.925 0.165 891.185 8.825 ;
      RECT 889.905 0.3 890.165 4.63 ;
      RECT 890.415 617.545 890.615 618.275 ;
      RECT 890.915 617.545 891.115 618.275 ;
      RECT 891.41 617.545 891.61 618.275 ;
      RECT 892.23 617.545 892.43 618.275 ;
      RECT 892.725 617.545 892.925 618.275 ;
      RECT 893.225 617.545 893.425 618.275 ;
      RECT 893.63 0.52 893.89 4.5 ;
      RECT 893.725 617.545 893.925 618.275 ;
      RECT 894.22 617.545 894.42 618.275 ;
      RECT 894.565 0.52 894.825 10.655 ;
      RECT 895.04 617.545 895.24 618.275 ;
      RECT 895.535 617.545 895.735 618.275 ;
      RECT 895.57 0.3 895.83 4.63 ;
      RECT 896.035 617.545 896.235 618.275 ;
      RECT 896.59 0.16 897.36 0.42 ;
      RECT 896.59 0.16 896.85 8.82 ;
      RECT 897.1 0.16 897.36 8.82 ;
      RECT 896.08 0.3 896.34 4.63 ;
      RECT 896.535 617.545 896.735 618.275 ;
      RECT 897.03 617.545 897.23 618.275 ;
      RECT 897.85 617.545 898.05 618.275 ;
      RECT 898.345 617.545 898.545 618.275 ;
      RECT 898.845 617.545 899.045 618.275 ;
      RECT 899.345 617.545 899.545 618.275 ;
      RECT 899.84 617.545 900.04 618.275 ;
      RECT 900.105 0.3 900.365 4.63 ;
      RECT 900.66 617.545 900.86 618.275 ;
      RECT 901.125 0.16 901.895 0.42 ;
      RECT 901.125 0.16 901.385 4.63 ;
      RECT 901.635 0.16 901.895 8.82 ;
      RECT 900.615 0.3 900.875 4.63 ;
      RECT 901.155 617.545 901.355 618.275 ;
      RECT 901.655 617.545 901.855 618.275 ;
      RECT 902.155 617.545 902.355 618.275 ;
      RECT 902.65 617.545 902.85 618.275 ;
      RECT 903.47 617.545 903.67 618.275 ;
      RECT 903.965 617.545 904.165 618.275 ;
      RECT 904.465 617.545 904.665 618.275 ;
      RECT 904.965 617.545 905.165 618.275 ;
      RECT 905.46 617.545 905.66 618.275 ;
      RECT 906.28 617.545 906.48 618.275 ;
      RECT 906.775 617.545 906.975 618.275 ;
      RECT 907.275 617.545 907.475 618.275 ;
      RECT 907.775 617.545 907.975 618.275 ;
      RECT 908.27 617.545 908.47 618.275 ;
      RECT 909.09 617.545 909.29 618.275 ;
      RECT 909.585 617.545 909.785 618.275 ;
      RECT 910.085 617.545 910.285 618.275 ;
      RECT 910.585 617.545 910.785 618.275 ;
      RECT 911.08 617.545 911.28 618.275 ;
      RECT 911.9 617.545 912.1 618.275 ;
      RECT 912.395 617.545 912.595 618.275 ;
      RECT 912.895 617.545 913.095 618.275 ;
      RECT 913.395 617.545 913.595 618.275 ;
      RECT 913.89 617.545 914.09 618.275 ;
      RECT 914.71 617.545 914.91 618.275 ;
      RECT 915.205 617.545 915.405 618.275 ;
      RECT 915.405 0.52 915.665 4.5 ;
      RECT 916.325 0.165 917.095 0.425 ;
      RECT 916.325 0.165 916.585 8.825 ;
      RECT 916.835 0.165 917.095 8.825 ;
      RECT 915.705 617.545 915.905 618.275 ;
      RECT 916.205 617.545 916.405 618.275 ;
      RECT 916.7 617.545 916.9 618.275 ;
      RECT 917.345 0.3 917.605 4.63 ;
      RECT 917.52 617.545 917.72 618.275 ;
      RECT 917.855 0.3 918.115 4.63 ;
      RECT 918.015 617.545 918.215 618.275 ;
      RECT 918.515 617.545 918.715 618.275 ;
      RECT 919.015 617.545 919.215 618.275 ;
      RECT 919.51 617.545 919.71 618.275 ;
      RECT 920.33 617.545 920.53 618.275 ;
      RECT 920.825 617.545 921.025 618.275 ;
      RECT 921.325 617.545 921.525 618.275 ;
      RECT 921.825 617.545 922.025 618.275 ;
      RECT 922.32 617.545 922.52 618.275 ;
      RECT 923.14 617.545 923.34 618.275 ;
      RECT 924.075 0.17 924.845 0.43 ;
      RECT 924.075 0.17 924.335 8.7 ;
      RECT 924.585 0.17 924.845 16.7 ;
      RECT 923.635 617.545 923.835 618.275 ;
      RECT 924.135 617.545 924.335 618.275 ;
      RECT 924.635 617.545 924.835 618.275 ;
      RECT 925.13 617.545 925.33 618.275 ;
      RECT 925.095 0.3 925.355 4.63 ;
      RECT 926.115 0.17 926.885 0.43 ;
      RECT 926.115 0.17 926.375 8.7 ;
      RECT 926.625 0.17 926.885 16.7 ;
      RECT 925.605 0.3 925.865 4.63 ;
      RECT 925.95 617.545 926.15 618.275 ;
      RECT 926.445 617.545 926.645 618.275 ;
      RECT 926.945 617.545 927.145 618.275 ;
      RECT 927.445 617.545 927.645 618.275 ;
      RECT 927.94 617.545 928.14 618.275 ;
      RECT 928.76 617.545 928.96 618.275 ;
      RECT 929.685 0.17 930.455 0.43 ;
      RECT 929.685 0.17 929.945 11.38 ;
      RECT 930.195 0.17 930.455 16.7 ;
      RECT 929.255 617.545 929.455 618.275 ;
      RECT 929.755 617.545 929.955 618.275 ;
      RECT 930.255 617.545 930.455 618.275 ;
      RECT 930.75 617.545 930.95 618.275 ;
      RECT 931.06 0.52 931.32 10.655 ;
      RECT 931.57 617.545 931.77 618.275 ;
      RECT 932.065 617.545 932.265 618.275 ;
      RECT 932.565 617.545 932.765 618.275 ;
      RECT 932.59 0.52 932.85 7.94 ;
      RECT 933.065 617.545 933.265 618.275 ;
      RECT 933.56 617.545 933.76 618.275 ;
      RECT 934.38 617.545 934.58 618.275 ;
      RECT 934.355 0.3 934.615 8.23 ;
      RECT 934.875 617.545 935.075 618.275 ;
      RECT 935.375 0.165 936.145 0.425 ;
      RECT 935.375 0.165 935.635 8.825 ;
      RECT 935.885 0.165 936.145 8.825 ;
      RECT 934.865 0.3 935.125 4.63 ;
      RECT 935.375 617.545 935.575 618.275 ;
      RECT 935.875 617.545 936.075 618.275 ;
      RECT 936.37 617.545 936.57 618.275 ;
      RECT 937.19 617.545 937.39 618.275 ;
      RECT 937.685 617.545 937.885 618.275 ;
      RECT 938.185 617.545 938.385 618.275 ;
      RECT 938.59 0.52 938.85 4.5 ;
      RECT 938.685 617.545 938.885 618.275 ;
      RECT 939.18 617.545 939.38 618.275 ;
      RECT 939.525 0.52 939.785 10.655 ;
      RECT 940 617.545 940.2 618.275 ;
      RECT 940.495 617.545 940.695 618.275 ;
      RECT 940.53 0.3 940.79 4.63 ;
      RECT 940.995 617.545 941.195 618.275 ;
      RECT 941.55 0.16 942.32 0.42 ;
      RECT 941.55 0.16 941.81 8.82 ;
      RECT 942.06 0.16 942.32 8.82 ;
      RECT 941.04 0.3 941.3 4.63 ;
      RECT 941.495 617.545 941.695 618.275 ;
      RECT 941.99 617.545 942.19 618.275 ;
      RECT 942.81 617.545 943.01 618.275 ;
      RECT 943.305 617.545 943.505 618.275 ;
      RECT 943.805 617.545 944.005 618.275 ;
      RECT 944.305 617.545 944.505 618.275 ;
      RECT 944.8 617.545 945 618.275 ;
      RECT 945.065 0.3 945.325 4.63 ;
      RECT 945.62 617.545 945.82 618.275 ;
      RECT 946.085 0.16 946.855 0.42 ;
      RECT 946.085 0.16 946.345 4.63 ;
      RECT 946.595 0.16 946.855 8.82 ;
      RECT 945.575 0.3 945.835 4.63 ;
      RECT 946.115 617.545 946.315 618.275 ;
      RECT 946.615 617.545 946.815 618.275 ;
      RECT 947.115 617.545 947.315 618.275 ;
      RECT 947.61 617.545 947.81 618.275 ;
      RECT 948.43 617.545 948.63 618.275 ;
      RECT 948.925 617.545 949.125 618.275 ;
      RECT 949.425 617.545 949.625 618.275 ;
      RECT 949.925 617.545 950.125 618.275 ;
      RECT 950.42 617.545 950.62 618.275 ;
      RECT 951.24 617.545 951.44 618.275 ;
      RECT 951.735 617.545 951.935 618.275 ;
      RECT 952.235 617.545 952.435 618.275 ;
      RECT 952.735 617.545 952.935 618.275 ;
      RECT 953.23 617.545 953.43 618.275 ;
      RECT 954.05 617.545 954.25 618.275 ;
      RECT 954.545 617.545 954.745 618.275 ;
      RECT 955.045 617.545 955.245 618.275 ;
      RECT 955.545 617.545 955.745 618.275 ;
      RECT 956.04 617.545 956.24 618.275 ;
      RECT 956.86 617.545 957.06 618.275 ;
      RECT 957.355 617.545 957.555 618.275 ;
      RECT 957.855 617.545 958.055 618.275 ;
      RECT 958.355 617.545 958.555 618.275 ;
      RECT 958.85 617.545 959.05 618.275 ;
      RECT 959.67 617.545 959.87 618.275 ;
      RECT 960.165 617.545 960.365 618.275 ;
      RECT 960.365 0.52 960.625 4.5 ;
      RECT 961.285 0.165 962.055 0.425 ;
      RECT 961.285 0.165 961.545 8.825 ;
      RECT 961.795 0.165 962.055 8.825 ;
      RECT 960.665 617.545 960.865 618.275 ;
      RECT 961.165 617.545 961.365 618.275 ;
      RECT 961.66 617.545 961.86 618.275 ;
      RECT 962.305 0.3 962.565 4.63 ;
      RECT 962.48 617.545 962.68 618.275 ;
      RECT 962.815 0.3 963.075 4.63 ;
      RECT 962.975 617.545 963.175 618.275 ;
      RECT 963.475 617.545 963.675 618.275 ;
      RECT 963.975 617.545 964.175 618.275 ;
      RECT 964.47 617.545 964.67 618.275 ;
      RECT 965.29 617.545 965.49 618.275 ;
      RECT 965.785 617.545 965.985 618.275 ;
      RECT 966.285 617.545 966.485 618.275 ;
      RECT 966.785 617.545 966.985 618.275 ;
      RECT 967.28 617.545 967.48 618.275 ;
      RECT 968.1 617.545 968.3 618.275 ;
      RECT 969.035 0.17 969.805 0.43 ;
      RECT 969.035 0.17 969.295 8.7 ;
      RECT 969.545 0.17 969.805 16.7 ;
      RECT 968.595 617.545 968.795 618.275 ;
      RECT 969.095 617.545 969.295 618.275 ;
      RECT 969.595 617.545 969.795 618.275 ;
      RECT 970.09 617.545 970.29 618.275 ;
      RECT 970.055 0.3 970.315 4.63 ;
      RECT 971.075 0.17 971.845 0.43 ;
      RECT 971.075 0.17 971.335 8.7 ;
      RECT 971.585 0.17 971.845 16.7 ;
      RECT 970.565 0.3 970.825 4.63 ;
      RECT 970.91 617.545 971.11 618.275 ;
      RECT 971.405 617.545 971.605 618.275 ;
      RECT 971.905 617.545 972.105 618.275 ;
      RECT 972.405 617.545 972.605 618.275 ;
      RECT 972.9 617.545 973.1 618.275 ;
      RECT 973.72 617.545 973.92 618.275 ;
      RECT 974.645 0.17 975.415 0.43 ;
      RECT 974.645 0.17 974.905 11.38 ;
      RECT 975.155 0.17 975.415 16.7 ;
      RECT 974.215 617.545 974.415 618.275 ;
      RECT 974.715 617.545 974.915 618.275 ;
      RECT 975.215 617.545 975.415 618.275 ;
      RECT 975.71 617.545 975.91 618.275 ;
      RECT 976.02 0.52 976.28 10.655 ;
      RECT 976.53 617.545 976.73 618.275 ;
      RECT 977.025 617.545 977.225 618.275 ;
      RECT 977.525 617.545 977.725 618.275 ;
      RECT 977.55 0.52 977.81 7.94 ;
      RECT 978.025 617.545 978.225 618.275 ;
      RECT 978.52 617.545 978.72 618.275 ;
      RECT 979.34 617.545 979.54 618.275 ;
      RECT 979.315 0.3 979.575 8.23 ;
      RECT 979.835 617.545 980.035 618.275 ;
      RECT 980.335 0.165 981.105 0.425 ;
      RECT 980.335 0.165 980.595 8.825 ;
      RECT 980.845 0.165 981.105 8.825 ;
      RECT 979.825 0.3 980.085 4.63 ;
      RECT 980.335 617.545 980.535 618.275 ;
      RECT 980.835 617.545 981.035 618.275 ;
      RECT 981.33 617.545 981.53 618.275 ;
      RECT 982.15 617.545 982.35 618.275 ;
      RECT 982.645 617.545 982.845 618.275 ;
      RECT 983.145 617.545 983.345 618.275 ;
      RECT 983.55 0.52 983.81 4.5 ;
      RECT 983.645 617.545 983.845 618.275 ;
      RECT 984.14 617.545 984.34 618.275 ;
      RECT 984.485 0.52 984.745 10.655 ;
      RECT 984.96 617.545 985.16 618.275 ;
      RECT 985.455 617.545 985.655 618.275 ;
      RECT 985.49 0.3 985.75 4.63 ;
      RECT 985.955 617.545 986.155 618.275 ;
      RECT 986.51 0.16 987.28 0.42 ;
      RECT 986.51 0.16 986.77 8.82 ;
      RECT 987.02 0.16 987.28 8.82 ;
      RECT 986 0.3 986.26 4.63 ;
      RECT 986.455 617.545 986.655 618.275 ;
      RECT 986.95 617.545 987.15 618.275 ;
      RECT 987.77 617.545 987.97 618.275 ;
      RECT 988.265 617.545 988.465 618.275 ;
      RECT 988.765 617.545 988.965 618.275 ;
      RECT 989.265 617.545 989.465 618.275 ;
      RECT 989.76 617.545 989.96 618.275 ;
      RECT 990.025 0.3 990.285 4.63 ;
      RECT 990.58 617.545 990.78 618.275 ;
      RECT 991.045 0.16 991.815 0.42 ;
      RECT 991.045 0.16 991.305 4.63 ;
      RECT 991.555 0.16 991.815 8.82 ;
      RECT 990.535 0.3 990.795 4.63 ;
      RECT 991.075 617.545 991.275 618.275 ;
      RECT 991.575 617.545 991.775 618.275 ;
      RECT 992.075 617.545 992.275 618.275 ;
      RECT 992.57 617.545 992.77 618.275 ;
      RECT 993.39 617.545 993.59 618.275 ;
      RECT 993.885 617.545 994.085 618.275 ;
      RECT 994.385 617.545 994.585 618.275 ;
      RECT 994.885 617.545 995.085 618.275 ;
      RECT 995.38 617.545 995.58 618.275 ;
      RECT 996.2 617.545 996.4 618.275 ;
      RECT 996.695 617.545 996.895 618.275 ;
      RECT 997.195 617.545 997.395 618.275 ;
      RECT 997.695 617.545 997.895 618.275 ;
      RECT 998.19 617.545 998.39 618.275 ;
      RECT 999.01 617.545 999.21 618.275 ;
      RECT 999.505 617.545 999.705 618.275 ;
      RECT 1000.005 617.545 1000.205 618.275 ;
      RECT 1000.505 617.545 1000.705 618.275 ;
      RECT 1001 617.545 1001.2 618.275 ;
      RECT 1001.82 617.545 1002.02 618.275 ;
      RECT 1002.315 617.545 1002.515 618.275 ;
      RECT 1002.815 617.545 1003.015 618.275 ;
      RECT 1003.315 617.545 1003.515 618.275 ;
      RECT 1003.81 617.545 1004.01 618.275 ;
      RECT 1004.63 617.545 1004.83 618.275 ;
      RECT 1005.125 617.545 1005.325 618.275 ;
      RECT 1005.325 0.52 1005.585 4.5 ;
      RECT 1006.245 0.165 1007.015 0.425 ;
      RECT 1006.245 0.165 1006.505 8.825 ;
      RECT 1006.755 0.165 1007.015 8.825 ;
      RECT 1005.625 617.545 1005.825 618.275 ;
      RECT 1006.125 617.545 1006.325 618.275 ;
      RECT 1006.62 617.545 1006.82 618.275 ;
      RECT 1007.265 0.3 1007.525 4.63 ;
      RECT 1007.44 617.545 1007.64 618.275 ;
      RECT 1007.775 0.3 1008.035 4.63 ;
      RECT 1007.935 617.545 1008.135 618.275 ;
      RECT 1008.435 617.545 1008.635 618.275 ;
      RECT 1008.935 617.545 1009.135 618.275 ;
      RECT 1009.43 617.545 1009.63 618.275 ;
      RECT 1010.25 617.545 1010.45 618.275 ;
      RECT 1010.745 617.545 1010.945 618.275 ;
      RECT 1011.245 617.545 1011.445 618.275 ;
      RECT 1011.745 617.545 1011.945 618.275 ;
      RECT 1012.24 617.545 1012.44 618.275 ;
      RECT 1013.06 617.545 1013.26 618.275 ;
      RECT 1013.995 0.17 1014.765 0.43 ;
      RECT 1013.995 0.17 1014.255 8.7 ;
      RECT 1014.505 0.17 1014.765 16.7 ;
      RECT 1013.555 617.545 1013.755 618.275 ;
      RECT 1014.055 617.545 1014.255 618.275 ;
      RECT 1014.555 617.545 1014.755 618.275 ;
      RECT 1015.05 617.545 1015.25 618.275 ;
      RECT 1015.015 0.3 1015.275 4.63 ;
      RECT 1016.035 0.17 1016.805 0.43 ;
      RECT 1016.035 0.17 1016.295 8.7 ;
      RECT 1016.545 0.17 1016.805 16.7 ;
      RECT 1015.525 0.3 1015.785 4.63 ;
      RECT 1015.87 617.545 1016.07 618.275 ;
      RECT 1016.365 617.545 1016.565 618.275 ;
      RECT 1016.865 617.545 1017.065 618.275 ;
      RECT 1017.365 617.545 1017.565 618.275 ;
      RECT 1017.86 617.545 1018.06 618.275 ;
      RECT 1018.68 617.545 1018.88 618.275 ;
      RECT 1019.605 0.17 1020.375 0.43 ;
      RECT 1019.605 0.17 1019.865 11.38 ;
      RECT 1020.115 0.17 1020.375 16.7 ;
      RECT 1019.175 617.545 1019.375 618.275 ;
      RECT 1019.675 617.545 1019.875 618.275 ;
      RECT 1020.175 617.545 1020.375 618.275 ;
      RECT 1020.67 617.545 1020.87 618.275 ;
      RECT 1020.98 0.52 1021.24 10.655 ;
      RECT 1021.49 617.545 1021.69 618.275 ;
      RECT 1021.985 617.545 1022.185 618.275 ;
      RECT 1022.485 617.545 1022.685 618.275 ;
      RECT 1022.51 0.52 1022.77 7.94 ;
      RECT 1022.985 617.545 1023.185 618.275 ;
      RECT 1023.48 617.545 1023.68 618.275 ;
      RECT 1024.3 617.545 1024.5 618.275 ;
      RECT 1024.275 0.3 1024.535 8.23 ;
      RECT 1024.795 617.545 1024.995 618.275 ;
      RECT 1025.295 0.165 1026.065 0.425 ;
      RECT 1025.295 0.165 1025.555 8.825 ;
      RECT 1025.805 0.165 1026.065 8.825 ;
      RECT 1024.785 0.3 1025.045 4.63 ;
      RECT 1025.295 617.545 1025.495 618.275 ;
      RECT 1025.795 617.545 1025.995 618.275 ;
      RECT 1026.29 617.545 1026.49 618.275 ;
      RECT 1027.11 617.545 1027.31 618.275 ;
      RECT 1027.605 617.545 1027.805 618.275 ;
      RECT 1028.105 617.545 1028.305 618.275 ;
      RECT 1028.51 0.52 1028.77 4.5 ;
      RECT 1028.605 617.545 1028.805 618.275 ;
      RECT 1029.1 617.545 1029.3 618.275 ;
      RECT 1029.445 0.52 1029.705 10.655 ;
      RECT 1029.92 617.545 1030.12 618.275 ;
      RECT 1030.415 617.545 1030.615 618.275 ;
      RECT 1030.45 0.3 1030.71 4.63 ;
      RECT 1030.915 617.545 1031.115 618.275 ;
      RECT 1031.47 0.16 1032.24 0.42 ;
      RECT 1031.47 0.16 1031.73 8.82 ;
      RECT 1031.98 0.16 1032.24 8.82 ;
      RECT 1030.96 0.3 1031.22 4.63 ;
      RECT 1031.415 617.545 1031.615 618.275 ;
      RECT 1031.91 617.545 1032.11 618.275 ;
      RECT 1032.73 617.545 1032.93 618.275 ;
      RECT 1033.225 617.545 1033.425 618.275 ;
      RECT 1033.725 617.545 1033.925 618.275 ;
      RECT 1034.225 617.545 1034.425 618.275 ;
      RECT 1034.72 617.545 1034.92 618.275 ;
      RECT 1034.985 0.3 1035.245 4.63 ;
      RECT 1035.54 617.545 1035.74 618.275 ;
      RECT 1036.005 0.16 1036.775 0.42 ;
      RECT 1036.005 0.16 1036.265 4.63 ;
      RECT 1036.515 0.16 1036.775 8.82 ;
      RECT 1035.495 0.3 1035.755 4.63 ;
      RECT 1036.035 617.545 1036.235 618.275 ;
      RECT 1036.535 617.545 1036.735 618.275 ;
      RECT 1037.035 617.545 1037.235 618.275 ;
      RECT 1037.53 617.545 1037.73 618.275 ;
      RECT 1038.35 617.545 1038.55 618.275 ;
      RECT 1038.845 617.545 1039.045 618.275 ;
      RECT 1039.345 617.545 1039.545 618.275 ;
      RECT 1039.845 617.545 1040.045 618.275 ;
      RECT 1040.34 617.545 1040.54 618.275 ;
      RECT 1041.16 617.545 1041.36 618.275 ;
      RECT 1041.655 617.545 1041.855 618.275 ;
      RECT 1042.155 617.545 1042.355 618.275 ;
      RECT 1042.655 617.545 1042.855 618.275 ;
      RECT 1043.15 617.545 1043.35 618.275 ;
      RECT 1043.97 617.545 1044.17 618.275 ;
      RECT 1044.465 617.545 1044.665 618.275 ;
      RECT 1044.965 617.545 1045.165 618.275 ;
      RECT 1045.465 617.545 1045.665 618.275 ;
      RECT 1045.96 617.545 1046.16 618.275 ;
      RECT 1046.78 617.545 1046.98 618.275 ;
      RECT 1047.275 617.545 1047.475 618.275 ;
      RECT 1047.775 617.545 1047.975 618.275 ;
      RECT 1048.275 617.545 1048.475 618.275 ;
      RECT 1048.77 617.545 1048.97 618.275 ;
      RECT 1049.59 617.545 1049.79 618.275 ;
      RECT 1050.085 617.545 1050.285 618.275 ;
      RECT 1050.285 0.52 1050.545 4.5 ;
      RECT 1051.205 0.165 1051.975 0.425 ;
      RECT 1051.205 0.165 1051.465 8.825 ;
      RECT 1051.715 0.165 1051.975 8.825 ;
      RECT 1050.585 617.545 1050.785 618.275 ;
      RECT 1051.085 617.545 1051.285 618.275 ;
      RECT 1051.58 617.545 1051.78 618.275 ;
      RECT 1052.225 0.3 1052.485 4.63 ;
      RECT 1052.4 617.545 1052.6 618.275 ;
      RECT 1052.735 0.3 1052.995 4.63 ;
      RECT 1052.895 617.545 1053.095 618.275 ;
      RECT 1053.395 617.545 1053.595 618.275 ;
      RECT 1053.895 617.545 1054.095 618.275 ;
      RECT 1054.39 617.545 1054.59 618.275 ;
      RECT 1055.21 617.545 1055.41 618.275 ;
      RECT 1055.705 617.545 1055.905 618.275 ;
      RECT 1056.205 617.545 1056.405 618.275 ;
      RECT 1056.705 617.545 1056.905 618.275 ;
      RECT 1057.2 617.545 1057.4 618.275 ;
      RECT 1058.02 617.545 1058.22 618.275 ;
      RECT 1058.955 0.17 1059.725 0.43 ;
      RECT 1058.955 0.17 1059.215 8.7 ;
      RECT 1059.465 0.17 1059.725 16.7 ;
      RECT 1058.515 617.545 1058.715 618.275 ;
      RECT 1059.015 617.545 1059.215 618.275 ;
      RECT 1059.515 617.545 1059.715 618.275 ;
      RECT 1060.01 617.545 1060.21 618.275 ;
      RECT 1059.975 0.3 1060.235 4.63 ;
      RECT 1060.995 0.17 1061.765 0.43 ;
      RECT 1060.995 0.17 1061.255 8.7 ;
      RECT 1061.505 0.17 1061.765 16.7 ;
      RECT 1060.485 0.3 1060.745 4.63 ;
      RECT 1060.83 617.545 1061.03 618.275 ;
      RECT 1061.325 617.545 1061.525 618.275 ;
      RECT 1061.825 617.545 1062.025 618.275 ;
      RECT 1062.325 617.545 1062.525 618.275 ;
      RECT 1062.82 617.545 1063.02 618.275 ;
      RECT 1063.64 617.545 1063.84 618.275 ;
      RECT 1064.565 0.17 1065.335 0.43 ;
      RECT 1064.565 0.17 1064.825 11.38 ;
      RECT 1065.075 0.17 1065.335 16.7 ;
      RECT 1064.135 617.545 1064.335 618.275 ;
      RECT 1064.635 617.545 1064.835 618.275 ;
      RECT 1065.135 617.545 1065.335 618.275 ;
      RECT 1065.63 617.545 1065.83 618.275 ;
      RECT 1065.94 0.52 1066.2 10.655 ;
      RECT 1066.45 617.545 1066.65 618.275 ;
      RECT 1066.945 617.545 1067.145 618.275 ;
      RECT 1067.445 617.545 1067.645 618.275 ;
      RECT 1067.47 0.52 1067.73 7.94 ;
      RECT 1067.945 617.545 1068.145 618.275 ;
      RECT 1068.44 617.545 1068.64 618.275 ;
      RECT 1069.26 617.545 1069.46 618.275 ;
      RECT 1069.235 0.3 1069.495 8.23 ;
      RECT 1069.755 617.545 1069.955 618.275 ;
      RECT 1070.255 0.165 1071.025 0.425 ;
      RECT 1070.255 0.165 1070.515 8.825 ;
      RECT 1070.765 0.165 1071.025 8.825 ;
      RECT 1069.745 0.3 1070.005 4.63 ;
      RECT 1070.255 617.545 1070.455 618.275 ;
      RECT 1070.755 617.545 1070.955 618.275 ;
      RECT 1071.25 617.545 1071.45 618.275 ;
      RECT 1072.07 617.545 1072.27 618.275 ;
      RECT 1072.565 617.545 1072.765 618.275 ;
      RECT 1073.065 617.545 1073.265 618.275 ;
      RECT 1073.47 0.52 1073.73 4.5 ;
      RECT 1073.565 617.545 1073.765 618.275 ;
      RECT 1074.06 617.545 1074.26 618.275 ;
      RECT 1074.405 0.52 1074.665 10.655 ;
      RECT 1074.88 617.545 1075.08 618.275 ;
      RECT 1075.375 617.545 1075.575 618.275 ;
      RECT 1075.41 0.3 1075.67 4.63 ;
      RECT 1075.875 617.545 1076.075 618.275 ;
      RECT 1076.43 0.16 1077.2 0.42 ;
      RECT 1076.43 0.16 1076.69 8.82 ;
      RECT 1076.94 0.16 1077.2 8.82 ;
      RECT 1075.92 0.3 1076.18 4.63 ;
      RECT 1076.375 617.545 1076.575 618.275 ;
      RECT 1076.87 617.545 1077.07 618.275 ;
      RECT 1077.69 617.545 1077.89 618.275 ;
      RECT 1078.185 617.545 1078.385 618.275 ;
      RECT 1078.685 617.545 1078.885 618.275 ;
      RECT 1079.185 617.545 1079.385 618.275 ;
      RECT 1079.68 617.545 1079.88 618.275 ;
      RECT 1079.945 0.3 1080.205 4.63 ;
      RECT 1080.5 617.545 1080.7 618.275 ;
      RECT 1080.965 0.16 1081.735 0.42 ;
      RECT 1080.965 0.16 1081.225 4.63 ;
      RECT 1081.475 0.16 1081.735 8.82 ;
      RECT 1080.455 0.3 1080.715 4.63 ;
      RECT 1080.995 617.545 1081.195 618.275 ;
      RECT 1081.495 617.545 1081.695 618.275 ;
      RECT 1081.995 617.545 1082.195 618.275 ;
      RECT 1082.49 617.545 1082.69 618.275 ;
      RECT 1083.31 617.545 1083.51 618.275 ;
      RECT 1083.805 617.545 1084.005 618.275 ;
      RECT 1084.305 617.545 1084.505 618.275 ;
      RECT 1084.805 617.545 1085.005 618.275 ;
      RECT 1085.3 617.545 1085.5 618.275 ;
      RECT 1086.12 617.545 1086.32 618.275 ;
      RECT 1086.615 617.545 1086.815 618.275 ;
      RECT 1087.115 617.545 1087.315 618.275 ;
      RECT 1087.615 617.545 1087.815 618.275 ;
      RECT 1088.11 617.545 1088.31 618.275 ;
      RECT 1088.93 617.545 1089.13 618.275 ;
      RECT 1089.425 617.545 1089.625 618.275 ;
      RECT 1089.925 617.545 1090.125 618.275 ;
      RECT 1090.425 617.545 1090.625 618.275 ;
      RECT 1090.92 617.545 1091.12 618.275 ;
      RECT 1091.74 617.545 1091.94 618.275 ;
      RECT 1092.235 617.545 1092.435 618.275 ;
      RECT 1092.735 617.545 1092.935 618.275 ;
      RECT 1093.235 617.545 1093.435 618.275 ;
      RECT 1093.73 617.545 1093.93 618.275 ;
      RECT 1094.55 617.545 1094.75 618.275 ;
      RECT 1095.045 617.545 1095.245 618.275 ;
      RECT 1095.245 0.52 1095.505 4.5 ;
      RECT 1096.165 0.165 1096.935 0.425 ;
      RECT 1096.165 0.165 1096.425 8.825 ;
      RECT 1096.675 0.165 1096.935 8.825 ;
      RECT 1095.545 617.545 1095.745 618.275 ;
      RECT 1096.045 617.545 1096.245 618.275 ;
      RECT 1096.54 617.545 1096.74 618.275 ;
      RECT 1097.185 0.3 1097.445 4.63 ;
      RECT 1097.36 617.545 1097.56 618.275 ;
      RECT 1097.695 0.3 1097.955 4.63 ;
      RECT 1097.855 617.545 1098.055 618.275 ;
      RECT 1098.355 617.545 1098.555 618.275 ;
      RECT 1098.855 617.545 1099.055 618.275 ;
      RECT 1099.35 617.545 1099.55 618.275 ;
      RECT 1100.17 617.545 1100.37 618.275 ;
      RECT 1100.665 617.545 1100.865 618.275 ;
      RECT 1101.165 617.545 1101.365 618.275 ;
      RECT 1101.665 617.545 1101.865 618.275 ;
      RECT 1102.16 617.545 1102.36 618.275 ;
      RECT 1102.98 617.545 1103.18 618.275 ;
      RECT 1103.915 0.17 1104.685 0.43 ;
      RECT 1103.915 0.17 1104.175 8.7 ;
      RECT 1104.425 0.17 1104.685 16.7 ;
      RECT 1103.475 617.545 1103.675 618.275 ;
      RECT 1103.975 617.545 1104.175 618.275 ;
      RECT 1104.475 617.545 1104.675 618.275 ;
      RECT 1104.97 617.545 1105.17 618.275 ;
      RECT 1104.935 0.3 1105.195 4.63 ;
      RECT 1105.955 0.17 1106.725 0.43 ;
      RECT 1105.955 0.17 1106.215 8.7 ;
      RECT 1106.465 0.17 1106.725 16.7 ;
      RECT 1105.445 0.3 1105.705 4.63 ;
      RECT 1105.79 617.545 1105.99 618.275 ;
      RECT 1106.285 617.545 1106.485 618.275 ;
      RECT 1106.785 617.545 1106.985 618.275 ;
      RECT 1107.285 617.545 1107.485 618.275 ;
      RECT 1107.78 617.545 1107.98 618.275 ;
      RECT 1108.6 617.545 1108.8 618.275 ;
      RECT 1109.525 0.17 1110.295 0.43 ;
      RECT 1109.525 0.17 1109.785 11.38 ;
      RECT 1110.035 0.17 1110.295 16.7 ;
      RECT 1109.095 617.545 1109.295 618.275 ;
      RECT 1109.595 617.545 1109.795 618.275 ;
      RECT 1110.095 617.545 1110.295 618.275 ;
      RECT 1110.59 617.545 1110.79 618.275 ;
      RECT 1110.9 0.52 1111.16 10.655 ;
      RECT 1111.41 617.545 1111.61 618.275 ;
      RECT 1111.905 617.545 1112.105 618.275 ;
      RECT 1112.405 617.545 1112.605 618.275 ;
      RECT 1112.43 0.52 1112.69 7.94 ;
      RECT 1112.905 617.545 1113.105 618.275 ;
      RECT 1113.4 617.545 1113.6 618.275 ;
      RECT 1114.22 617.545 1114.42 618.275 ;
      RECT 1114.195 0.3 1114.455 8.23 ;
      RECT 1114.715 617.545 1114.915 618.275 ;
      RECT 1115.215 0.165 1115.985 0.425 ;
      RECT 1115.215 0.165 1115.475 8.825 ;
      RECT 1115.725 0.165 1115.985 8.825 ;
      RECT 1114.705 0.3 1114.965 4.63 ;
      RECT 1115.215 617.545 1115.415 618.275 ;
      RECT 1115.715 617.545 1115.915 618.275 ;
      RECT 1116.21 617.545 1116.41 618.275 ;
      RECT 1117.03 617.545 1117.23 618.275 ;
      RECT 1117.525 617.545 1117.725 618.275 ;
      RECT 1118.025 617.545 1118.225 618.275 ;
      RECT 1118.43 0.52 1118.69 4.5 ;
      RECT 1118.525 617.545 1118.725 618.275 ;
      RECT 1119.02 617.545 1119.22 618.275 ;
      RECT 1119.365 0.52 1119.625 10.655 ;
      RECT 1119.84 617.545 1120.04 618.275 ;
      RECT 1120.335 617.545 1120.535 618.275 ;
      RECT 1120.37 0.3 1120.63 4.63 ;
      RECT 1120.835 617.545 1121.035 618.275 ;
      RECT 1121.39 0.16 1122.16 0.42 ;
      RECT 1121.39 0.16 1121.65 8.82 ;
      RECT 1121.9 0.16 1122.16 8.82 ;
      RECT 1120.88 0.3 1121.14 4.63 ;
      RECT 1121.335 617.545 1121.535 618.275 ;
      RECT 1121.83 617.545 1122.03 618.275 ;
      RECT 1122.65 617.545 1122.85 618.275 ;
      RECT 1123.145 617.545 1123.345 618.275 ;
      RECT 1123.645 617.545 1123.845 618.275 ;
      RECT 1124.145 617.545 1124.345 618.275 ;
      RECT 1124.64 617.545 1124.84 618.275 ;
      RECT 1124.905 0.3 1125.165 4.63 ;
      RECT 1125.46 617.545 1125.66 618.275 ;
      RECT 1125.925 0.16 1126.695 0.42 ;
      RECT 1125.925 0.16 1126.185 4.63 ;
      RECT 1126.435 0.16 1126.695 8.82 ;
      RECT 1125.415 0.3 1125.675 4.63 ;
      RECT 1125.955 617.545 1126.155 618.275 ;
      RECT 1126.455 617.545 1126.655 618.275 ;
      RECT 1126.955 617.545 1127.155 618.275 ;
      RECT 1127.45 617.545 1127.65 618.275 ;
      RECT 1128.27 617.545 1128.47 618.275 ;
      RECT 1128.765 617.545 1128.965 618.275 ;
      RECT 1129.265 617.545 1129.465 618.275 ;
      RECT 1129.765 617.545 1129.965 618.275 ;
      RECT 1130.26 617.545 1130.46 618.275 ;
      RECT 1131.08 617.545 1131.28 618.275 ;
      RECT 1131.575 617.545 1131.775 618.275 ;
      RECT 1132.075 617.545 1132.275 618.275 ;
      RECT 1132.575 617.545 1132.775 618.275 ;
      RECT 1133.07 617.545 1133.27 618.275 ;
      RECT 1133.89 617.545 1134.09 618.275 ;
      RECT 1134.385 617.545 1134.585 618.275 ;
      RECT 1134.885 617.545 1135.085 618.275 ;
      RECT 1135.385 617.545 1135.585 618.275 ;
      RECT 1135.88 617.545 1136.08 618.275 ;
      RECT 1136.7 617.545 1136.9 618.275 ;
      RECT 1137.195 617.545 1137.395 618.275 ;
      RECT 1137.695 617.545 1137.895 618.275 ;
      RECT 1138.195 617.545 1138.395 618.275 ;
      RECT 1138.69 617.545 1138.89 618.275 ;
      RECT 1139.51 617.545 1139.71 618.275 ;
      RECT 1140.005 617.545 1140.205 618.275 ;
      RECT 1140.205 0.52 1140.465 4.5 ;
      RECT 1141.125 0.165 1141.895 0.425 ;
      RECT 1141.125 0.165 1141.385 8.825 ;
      RECT 1141.635 0.165 1141.895 8.825 ;
      RECT 1140.505 617.545 1140.705 618.275 ;
      RECT 1141.005 617.545 1141.205 618.275 ;
      RECT 1141.5 617.545 1141.7 618.275 ;
      RECT 1142.145 0.3 1142.405 4.63 ;
      RECT 1142.32 617.545 1142.52 618.275 ;
      RECT 1142.655 0.3 1142.915 4.63 ;
      RECT 1142.815 617.545 1143.015 618.275 ;
      RECT 1143.315 617.545 1143.515 618.275 ;
      RECT 1143.815 617.545 1144.015 618.275 ;
      RECT 1144.31 617.545 1144.51 618.275 ;
      RECT 1145.13 617.545 1145.33 618.275 ;
      RECT 1145.625 617.545 1145.825 618.275 ;
      RECT 1146.125 617.545 1146.325 618.275 ;
      RECT 1146.625 617.545 1146.825 618.275 ;
      RECT 1147.12 617.545 1147.32 618.275 ;
      RECT 1147.94 617.545 1148.14 618.275 ;
      RECT 1148.875 0.17 1149.645 0.43 ;
      RECT 1148.875 0.17 1149.135 8.7 ;
      RECT 1149.385 0.17 1149.645 16.7 ;
      RECT 1148.435 617.545 1148.635 618.275 ;
      RECT 1148.935 617.545 1149.135 618.275 ;
      RECT 1149.435 617.545 1149.635 618.275 ;
      RECT 1149.93 617.545 1150.13 618.275 ;
      RECT 1149.895 0.3 1150.155 4.63 ;
      RECT 1150.915 0.17 1151.685 0.43 ;
      RECT 1150.915 0.17 1151.175 8.7 ;
      RECT 1151.425 0.17 1151.685 16.7 ;
      RECT 1150.405 0.3 1150.665 4.63 ;
      RECT 1150.75 617.545 1150.95 618.275 ;
      RECT 1151.245 617.545 1151.445 618.275 ;
      RECT 1151.745 617.545 1151.945 618.275 ;
      RECT 1152.245 617.545 1152.445 618.275 ;
      RECT 1152.74 617.545 1152.94 618.275 ;
      RECT 1153.56 617.545 1153.76 618.275 ;
      RECT 1154.485 0.17 1155.255 0.43 ;
      RECT 1154.485 0.17 1154.745 11.38 ;
      RECT 1154.995 0.17 1155.255 16.7 ;
      RECT 1154.055 617.545 1154.255 618.275 ;
      RECT 1154.555 617.545 1154.755 618.275 ;
      RECT 1155.055 617.545 1155.255 618.275 ;
      RECT 1155.55 617.545 1155.75 618.275 ;
      RECT 1155.86 0.52 1156.12 10.655 ;
      RECT 1156.37 617.545 1156.57 618.275 ;
      RECT 1156.865 617.545 1157.065 618.275 ;
      RECT 1157.365 617.545 1157.565 618.275 ;
      RECT 1157.39 0.52 1157.65 7.94 ;
      RECT 1157.865 617.545 1158.065 618.275 ;
      RECT 1158.36 617.545 1158.56 618.275 ;
      RECT 1159.18 617.545 1159.38 618.275 ;
      RECT 1159.155 0.3 1159.415 8.23 ;
      RECT 1159.675 617.545 1159.875 618.275 ;
      RECT 1160.175 0.165 1160.945 0.425 ;
      RECT 1160.175 0.165 1160.435 8.825 ;
      RECT 1160.685 0.165 1160.945 8.825 ;
      RECT 1159.665 0.3 1159.925 4.63 ;
      RECT 1160.175 617.545 1160.375 618.275 ;
      RECT 1160.675 617.545 1160.875 618.275 ;
      RECT 1161.17 617.545 1161.37 618.275 ;
      RECT 1161.99 617.545 1162.19 618.275 ;
      RECT 1162.485 617.545 1162.685 618.275 ;
      RECT 1162.985 617.545 1163.185 618.275 ;
      RECT 1163.39 0.52 1163.65 4.5 ;
      RECT 1163.485 617.545 1163.685 618.275 ;
      RECT 1163.98 617.545 1164.18 618.275 ;
      RECT 1164.325 0.52 1164.585 10.655 ;
      RECT 1164.8 617.545 1165 618.275 ;
      RECT 1165.295 617.545 1165.495 618.275 ;
      RECT 1165.33 0.3 1165.59 4.63 ;
      RECT 1165.795 617.545 1165.995 618.275 ;
      RECT 1166.35 0.16 1167.12 0.42 ;
      RECT 1166.35 0.16 1166.61 8.82 ;
      RECT 1166.86 0.16 1167.12 8.82 ;
      RECT 1165.84 0.3 1166.1 4.63 ;
      RECT 1166.295 617.545 1166.495 618.275 ;
      RECT 1166.79 617.545 1166.99 618.275 ;
      RECT 1167.61 617.545 1167.81 618.275 ;
      RECT 1168.105 617.545 1168.305 618.275 ;
      RECT 1168.605 617.545 1168.805 618.275 ;
      RECT 1169.105 617.545 1169.305 618.275 ;
      RECT 1169.6 617.545 1169.8 618.275 ;
      RECT 1169.865 0.3 1170.125 4.63 ;
      RECT 1170.42 617.545 1170.62 618.275 ;
      RECT 1170.885 0.16 1171.655 0.42 ;
      RECT 1170.885 0.16 1171.145 4.63 ;
      RECT 1171.395 0.16 1171.655 8.82 ;
      RECT 1170.375 0.3 1170.635 4.63 ;
      RECT 1170.915 617.545 1171.115 618.275 ;
      RECT 1171.415 617.545 1171.615 618.275 ;
      RECT 1171.915 617.545 1172.115 618.275 ;
      RECT 1172.41 617.545 1172.61 618.275 ;
      RECT 1173.23 617.545 1173.43 618.275 ;
      RECT 1173.725 617.545 1173.925 618.275 ;
      RECT 1174.225 617.545 1174.425 618.275 ;
      RECT 1174.725 617.545 1174.925 618.275 ;
      RECT 1175.22 617.545 1175.42 618.275 ;
      RECT 1176.04 617.545 1176.24 618.275 ;
      RECT 1176.535 617.545 1176.735 618.275 ;
      RECT 1177.035 617.545 1177.235 618.275 ;
      RECT 1177.535 617.545 1177.735 618.275 ;
      RECT 1178.03 617.545 1178.23 618.275 ;
      RECT 1178.85 617.545 1179.05 618.275 ;
      RECT 1179.345 617.545 1179.545 618.275 ;
      RECT 1179.845 617.545 1180.045 618.275 ;
      RECT 1180.345 617.545 1180.545 618.275 ;
      RECT 1180.84 617.545 1181.04 618.275 ;
      RECT 1181.66 617.545 1181.86 618.275 ;
      RECT 1182.155 617.545 1182.355 618.275 ;
      RECT 1182.655 617.545 1182.855 618.275 ;
      RECT 1183.155 617.545 1183.355 618.275 ;
      RECT 1183.65 617.545 1183.85 618.275 ;
      RECT 1184.47 617.545 1184.67 618.275 ;
      RECT 1184.965 617.545 1185.165 618.275 ;
      RECT 1185.165 0.52 1185.425 4.5 ;
      RECT 1186.085 0.165 1186.855 0.425 ;
      RECT 1186.085 0.165 1186.345 8.825 ;
      RECT 1186.595 0.165 1186.855 8.825 ;
      RECT 1185.465 617.545 1185.665 618.275 ;
      RECT 1185.965 617.545 1186.165 618.275 ;
      RECT 1186.46 617.545 1186.66 618.275 ;
      RECT 1187.105 0.3 1187.365 4.63 ;
      RECT 1187.28 617.545 1187.48 618.275 ;
      RECT 1187.615 0.3 1187.875 4.63 ;
      RECT 1187.775 617.545 1187.975 618.275 ;
      RECT 1188.275 617.545 1188.475 618.275 ;
      RECT 1188.775 617.545 1188.975 618.275 ;
      RECT 1189.27 617.545 1189.47 618.275 ;
      RECT 1190.09 617.545 1190.29 618.275 ;
      RECT 1190.585 617.545 1190.785 618.275 ;
      RECT 1191.085 617.545 1191.285 618.275 ;
      RECT 1191.585 617.545 1191.785 618.275 ;
      RECT 1192.08 617.545 1192.28 618.275 ;
      RECT 1192.9 617.545 1193.1 618.275 ;
      RECT 1193.835 0.17 1194.605 0.43 ;
      RECT 1193.835 0.17 1194.095 8.7 ;
      RECT 1194.345 0.17 1194.605 16.7 ;
      RECT 1193.395 617.545 1193.595 618.275 ;
      RECT 1193.895 617.545 1194.095 618.275 ;
      RECT 1194.395 617.545 1194.595 618.275 ;
      RECT 1194.89 617.545 1195.09 618.275 ;
      RECT 1194.855 0.3 1195.115 4.63 ;
      RECT 1195.875 0.17 1196.645 0.43 ;
      RECT 1195.875 0.17 1196.135 8.7 ;
      RECT 1196.385 0.17 1196.645 16.7 ;
      RECT 1195.365 0.3 1195.625 4.63 ;
      RECT 1195.71 617.545 1195.91 618.275 ;
      RECT 1196.205 617.545 1196.405 618.275 ;
      RECT 1196.705 617.545 1196.905 618.275 ;
      RECT 1197.205 617.545 1197.405 618.275 ;
      RECT 1197.7 617.545 1197.9 618.275 ;
      RECT 1198.52 617.545 1198.72 618.275 ;
      RECT 1199.445 0.17 1200.215 0.43 ;
      RECT 1199.445 0.17 1199.705 11.38 ;
      RECT 1199.955 0.17 1200.215 16.7 ;
      RECT 1199.015 617.545 1199.215 618.275 ;
      RECT 1199.515 617.545 1199.715 618.275 ;
      RECT 1200.015 617.545 1200.215 618.275 ;
      RECT 1200.51 617.545 1200.71 618.275 ;
      RECT 1200.82 0.52 1201.08 10.655 ;
      RECT 1201.33 617.545 1201.53 618.275 ;
      RECT 1201.825 617.545 1202.025 618.275 ;
      RECT 1202.325 617.545 1202.525 618.275 ;
      RECT 1202.35 0.52 1202.61 7.94 ;
      RECT 1202.825 617.545 1203.025 618.275 ;
      RECT 1203.32 617.545 1203.52 618.275 ;
      RECT 1204.14 617.545 1204.34 618.275 ;
      RECT 1204.115 0.3 1204.375 8.23 ;
      RECT 1204.635 617.545 1204.835 618.275 ;
      RECT 1205.135 0.165 1205.905 0.425 ;
      RECT 1205.135 0.165 1205.395 8.825 ;
      RECT 1205.645 0.165 1205.905 8.825 ;
      RECT 1204.625 0.3 1204.885 4.63 ;
      RECT 1205.135 617.545 1205.335 618.275 ;
      RECT 1205.635 617.545 1205.835 618.275 ;
      RECT 1206.13 617.545 1206.33 618.275 ;
      RECT 1206.95 617.545 1207.15 618.275 ;
      RECT 1207.445 617.545 1207.645 618.275 ;
      RECT 1207.945 617.545 1208.145 618.275 ;
      RECT 1208.35 0.52 1208.61 4.5 ;
      RECT 1208.445 617.545 1208.645 618.275 ;
      RECT 1208.94 617.545 1209.14 618.275 ;
      RECT 1209.285 0.52 1209.545 10.655 ;
      RECT 1209.76 617.545 1209.96 618.275 ;
      RECT 1210.255 617.545 1210.455 618.275 ;
      RECT 1210.29 0.3 1210.55 4.63 ;
      RECT 1210.755 617.545 1210.955 618.275 ;
      RECT 1211.31 0.16 1212.08 0.42 ;
      RECT 1211.31 0.16 1211.57 8.82 ;
      RECT 1211.82 0.16 1212.08 8.82 ;
      RECT 1210.8 0.3 1211.06 4.63 ;
      RECT 1211.255 617.545 1211.455 618.275 ;
      RECT 1211.75 617.545 1211.95 618.275 ;
      RECT 1212.57 617.545 1212.77 618.275 ;
      RECT 1213.065 617.545 1213.265 618.275 ;
      RECT 1213.565 617.545 1213.765 618.275 ;
      RECT 1214.065 617.545 1214.265 618.275 ;
      RECT 1214.56 617.545 1214.76 618.275 ;
      RECT 1214.825 0.3 1215.085 4.63 ;
      RECT 1215.38 617.545 1215.58 618.275 ;
      RECT 1215.845 0.16 1216.615 0.42 ;
      RECT 1215.845 0.16 1216.105 4.63 ;
      RECT 1216.355 0.16 1216.615 8.82 ;
      RECT 1215.335 0.3 1215.595 4.63 ;
      RECT 1215.875 617.545 1216.075 618.275 ;
      RECT 1216.375 617.545 1216.575 618.275 ;
      RECT 1216.875 617.545 1217.075 618.275 ;
      RECT 1217.37 617.545 1217.57 618.275 ;
      RECT 1218.19 617.545 1218.39 618.275 ;
      RECT 1218.685 617.545 1218.885 618.275 ;
      RECT 1219.185 617.545 1219.385 618.275 ;
      RECT 1219.685 617.545 1219.885 618.275 ;
      RECT 1220.18 617.545 1220.38 618.275 ;
      RECT 1221 617.545 1221.2 618.275 ;
      RECT 1221.495 617.545 1221.695 618.275 ;
      RECT 1221.995 617.545 1222.195 618.275 ;
      RECT 1222.495 617.545 1222.695 618.275 ;
      RECT 1222.99 617.545 1223.19 618.275 ;
      RECT 1223.81 617.545 1224.01 618.275 ;
      RECT 1224.305 617.545 1224.505 618.275 ;
      RECT 1224.805 617.545 1225.005 618.275 ;
      RECT 1225.305 617.545 1225.505 618.275 ;
      RECT 1225.8 617.545 1226 618.275 ;
      RECT 1226.62 617.545 1226.82 618.275 ;
      RECT 1227.115 617.545 1227.315 618.275 ;
      RECT 1227.615 617.545 1227.815 618.275 ;
      RECT 1228.115 617.545 1228.315 618.275 ;
      RECT 1228.61 617.545 1228.81 618.275 ;
      RECT 1229.43 617.545 1229.63 618.275 ;
      RECT 1229.925 617.545 1230.125 618.275 ;
      RECT 1230.125 0.52 1230.385 4.5 ;
      RECT 1231.045 0.165 1231.815 0.425 ;
      RECT 1231.045 0.165 1231.305 8.825 ;
      RECT 1231.555 0.165 1231.815 8.825 ;
      RECT 1230.425 617.545 1230.625 618.275 ;
      RECT 1230.925 617.545 1231.125 618.275 ;
      RECT 1231.42 617.545 1231.62 618.275 ;
      RECT 1232.065 0.3 1232.325 4.63 ;
      RECT 1232.24 617.545 1232.44 618.275 ;
      RECT 1232.575 0.3 1232.835 4.63 ;
      RECT 1232.735 617.545 1232.935 618.275 ;
      RECT 1233.235 617.545 1233.435 618.275 ;
      RECT 1233.735 617.545 1233.935 618.275 ;
      RECT 1234.23 617.545 1234.43 618.275 ;
      RECT 1235.05 617.545 1235.25 618.275 ;
      RECT 1235.545 617.545 1235.745 618.275 ;
      RECT 1236.045 617.545 1236.245 618.275 ;
      RECT 1236.545 617.545 1236.745 618.275 ;
      RECT 1237.04 617.545 1237.24 618.275 ;
      RECT 1237.86 617.545 1238.06 618.275 ;
      RECT 1238.795 0.17 1239.565 0.43 ;
      RECT 1238.795 0.17 1239.055 8.7 ;
      RECT 1239.305 0.17 1239.565 16.7 ;
      RECT 1238.355 617.545 1238.555 618.275 ;
      RECT 1238.855 617.545 1239.055 618.275 ;
      RECT 1239.355 617.545 1239.555 618.275 ;
      RECT 1239.85 617.545 1240.05 618.275 ;
      RECT 1239.815 0.3 1240.075 4.63 ;
      RECT 1240.835 0.17 1241.605 0.43 ;
      RECT 1240.835 0.17 1241.095 8.7 ;
      RECT 1241.345 0.17 1241.605 16.7 ;
      RECT 1240.325 0.3 1240.585 4.63 ;
      RECT 1240.67 617.545 1240.87 618.275 ;
      RECT 1241.165 617.545 1241.365 618.275 ;
      RECT 1241.665 617.545 1241.865 618.275 ;
      RECT 1242.165 617.545 1242.365 618.275 ;
      RECT 1242.66 617.545 1242.86 618.275 ;
      RECT 1243.48 617.545 1243.68 618.275 ;
      RECT 1244.405 0.17 1245.175 0.43 ;
      RECT 1244.405 0.17 1244.665 11.38 ;
      RECT 1244.915 0.17 1245.175 16.7 ;
      RECT 1243.975 617.545 1244.175 618.275 ;
      RECT 1244.475 617.545 1244.675 618.275 ;
      RECT 1244.975 617.545 1245.175 618.275 ;
      RECT 1245.47 617.545 1245.67 618.275 ;
      RECT 1245.78 0.52 1246.04 10.655 ;
      RECT 1246.29 617.545 1246.49 618.275 ;
      RECT 1246.785 617.545 1246.985 618.275 ;
      RECT 1247.285 617.545 1247.485 618.275 ;
      RECT 1247.31 0.52 1247.57 7.94 ;
      RECT 1247.785 617.545 1247.985 618.275 ;
      RECT 1248.28 617.545 1248.48 618.275 ;
      RECT 1249.1 617.545 1249.3 618.275 ;
      RECT 1249.075 0.3 1249.335 8.23 ;
      RECT 1249.595 617.545 1249.795 618.275 ;
      RECT 1250.095 0.165 1250.865 0.425 ;
      RECT 1250.095 0.165 1250.355 8.825 ;
      RECT 1250.605 0.165 1250.865 8.825 ;
      RECT 1249.585 0.3 1249.845 4.63 ;
      RECT 1250.095 617.545 1250.295 618.275 ;
      RECT 1250.595 617.545 1250.795 618.275 ;
      RECT 1251.09 617.545 1251.29 618.275 ;
      RECT 1251.91 617.545 1252.11 618.275 ;
      RECT 1252.405 617.545 1252.605 618.275 ;
      RECT 1252.905 617.545 1253.105 618.275 ;
      RECT 1253.31 0.52 1253.57 4.5 ;
      RECT 1253.405 617.545 1253.605 618.275 ;
      RECT 1253.9 617.545 1254.1 618.275 ;
      RECT 1254.245 0.52 1254.505 10.655 ;
      RECT 1254.72 617.545 1254.92 618.275 ;
      RECT 1255.215 617.545 1255.415 618.275 ;
      RECT 1255.25 0.3 1255.51 4.63 ;
      RECT 1255.715 617.545 1255.915 618.275 ;
      RECT 1256.27 0.16 1257.04 0.42 ;
      RECT 1256.27 0.16 1256.53 8.82 ;
      RECT 1256.78 0.16 1257.04 8.82 ;
      RECT 1255.76 0.3 1256.02 4.63 ;
      RECT 1256.215 617.545 1256.415 618.275 ;
      RECT 1256.71 617.545 1256.91 618.275 ;
      RECT 1257.53 617.545 1257.73 618.275 ;
      RECT 1258.025 617.545 1258.225 618.275 ;
      RECT 1258.525 617.545 1258.725 618.275 ;
      RECT 1259.025 617.545 1259.225 618.275 ;
      RECT 1259.52 617.545 1259.72 618.275 ;
      RECT 1259.785 0.3 1260.045 4.63 ;
      RECT 1260.34 617.545 1260.54 618.275 ;
      RECT 1260.805 0.16 1261.575 0.42 ;
      RECT 1260.805 0.16 1261.065 4.63 ;
      RECT 1261.315 0.16 1261.575 8.82 ;
      RECT 1260.295 0.3 1260.555 4.63 ;
      RECT 1260.835 617.545 1261.035 618.275 ;
      RECT 1261.335 617.545 1261.535 618.275 ;
      RECT 1261.835 617.545 1262.035 618.275 ;
      RECT 1262.33 617.545 1262.53 618.275 ;
      RECT 1263.15 617.545 1263.35 618.275 ;
      RECT 1263.645 617.545 1263.845 618.275 ;
      RECT 1264.145 617.545 1264.345 618.275 ;
      RECT 1264.645 617.545 1264.845 618.275 ;
      RECT 1265.14 617.545 1265.34 618.275 ;
      RECT 1265.96 617.545 1266.16 618.275 ;
      RECT 1266.455 617.545 1266.655 618.275 ;
      RECT 1266.955 617.545 1267.155 618.275 ;
      RECT 1267.455 617.545 1267.655 618.275 ;
      RECT 1267.95 617.545 1268.15 618.275 ;
      RECT 1268.77 617.545 1268.97 618.275 ;
      RECT 1269.265 617.545 1269.465 618.275 ;
      RECT 1269.765 617.545 1269.965 618.275 ;
      RECT 1270.265 617.545 1270.465 618.275 ;
      RECT 1270.76 617.545 1270.96 618.275 ;
      RECT 1271.58 617.545 1271.78 618.275 ;
      RECT 1272.075 617.545 1272.275 618.275 ;
      RECT 1272.575 617.545 1272.775 618.275 ;
      RECT 1273.075 617.545 1273.275 618.275 ;
      RECT 1273.57 617.545 1273.77 618.275 ;
      RECT 1274.39 617.545 1274.59 618.275 ;
      RECT 1274.885 617.545 1275.085 618.275 ;
      RECT 1275.085 0.52 1275.345 4.5 ;
      RECT 1276.005 0.165 1276.775 0.425 ;
      RECT 1276.005 0.165 1276.265 8.825 ;
      RECT 1276.515 0.165 1276.775 8.825 ;
      RECT 1275.385 617.545 1275.585 618.275 ;
      RECT 1275.885 617.545 1276.085 618.275 ;
      RECT 1276.38 617.545 1276.58 618.275 ;
      RECT 1277.025 0.3 1277.285 4.63 ;
      RECT 1277.2 617.545 1277.4 618.275 ;
      RECT 1277.535 0.3 1277.795 4.63 ;
      RECT 1277.695 617.545 1277.895 618.275 ;
      RECT 1278.195 617.545 1278.395 618.275 ;
      RECT 1278.695 617.545 1278.895 618.275 ;
      RECT 1279.19 617.545 1279.39 618.275 ;
      RECT 1280.01 617.545 1280.21 618.275 ;
      RECT 1280.505 617.545 1280.705 618.275 ;
      RECT 1281.005 617.545 1281.205 618.275 ;
      RECT 1281.505 617.545 1281.705 618.275 ;
      RECT 1282 617.545 1282.2 618.275 ;
      RECT 1282.82 617.545 1283.02 618.275 ;
      RECT 1283.755 0.17 1284.525 0.43 ;
      RECT 1283.755 0.17 1284.015 8.7 ;
      RECT 1284.265 0.17 1284.525 16.7 ;
      RECT 1283.315 617.545 1283.515 618.275 ;
      RECT 1283.815 617.545 1284.015 618.275 ;
      RECT 1284.315 617.545 1284.515 618.275 ;
      RECT 1284.81 617.545 1285.01 618.275 ;
      RECT 1284.775 0.3 1285.035 4.63 ;
      RECT 1285.795 0.17 1286.565 0.43 ;
      RECT 1285.795 0.17 1286.055 8.7 ;
      RECT 1286.305 0.17 1286.565 16.7 ;
      RECT 1285.285 0.3 1285.545 4.63 ;
      RECT 1285.63 617.545 1285.83 618.275 ;
      RECT 1286.125 617.545 1286.325 618.275 ;
      RECT 1286.625 617.545 1286.825 618.275 ;
      RECT 1287.125 617.545 1287.325 618.275 ;
      RECT 1287.62 617.545 1287.82 618.275 ;
      RECT 1288.44 617.545 1288.64 618.275 ;
      RECT 1289.365 0.17 1290.135 0.43 ;
      RECT 1289.365 0.17 1289.625 11.38 ;
      RECT 1289.875 0.17 1290.135 16.7 ;
      RECT 1288.935 617.545 1289.135 618.275 ;
      RECT 1289.435 617.545 1289.635 618.275 ;
      RECT 1289.935 617.545 1290.135 618.275 ;
      RECT 1290.43 617.545 1290.63 618.275 ;
      RECT 1290.74 0.52 1291 10.655 ;
      RECT 1291.25 617.545 1291.45 618.275 ;
      RECT 1291.745 617.545 1291.945 618.275 ;
      RECT 1292.245 617.545 1292.445 618.275 ;
      RECT 1292.27 0.52 1292.53 7.94 ;
      RECT 1292.745 617.545 1292.945 618.275 ;
      RECT 1293.24 617.545 1293.44 618.275 ;
      RECT 1294.06 617.545 1294.26 618.275 ;
      RECT 1294.035 0.3 1294.295 8.23 ;
      RECT 1294.555 617.545 1294.755 618.275 ;
      RECT 1295.055 0.165 1295.825 0.425 ;
      RECT 1295.055 0.165 1295.315 8.825 ;
      RECT 1295.565 0.165 1295.825 8.825 ;
      RECT 1294.545 0.3 1294.805 4.63 ;
      RECT 1295.055 617.545 1295.255 618.275 ;
      RECT 1295.555 617.545 1295.755 618.275 ;
      RECT 1296.05 617.545 1296.25 618.275 ;
      RECT 1296.87 617.545 1297.07 618.275 ;
      RECT 1297.365 617.545 1297.565 618.275 ;
      RECT 1297.865 617.545 1298.065 618.275 ;
      RECT 1298.27 0.52 1298.53 4.5 ;
      RECT 1298.365 617.545 1298.565 618.275 ;
      RECT 1298.86 617.545 1299.06 618.275 ;
      RECT 1299.205 0.52 1299.465 10.655 ;
      RECT 1299.68 617.545 1299.88 618.275 ;
      RECT 1300.175 617.545 1300.375 618.275 ;
      RECT 1300.21 0.3 1300.47 4.63 ;
      RECT 1300.675 617.545 1300.875 618.275 ;
      RECT 1301.23 0.16 1302 0.42 ;
      RECT 1301.23 0.16 1301.49 8.82 ;
      RECT 1301.74 0.16 1302 8.82 ;
      RECT 1300.72 0.3 1300.98 4.63 ;
      RECT 1301.175 617.545 1301.375 618.275 ;
      RECT 1301.67 617.545 1301.87 618.275 ;
      RECT 1302.49 617.545 1302.69 618.275 ;
      RECT 1302.985 617.545 1303.185 618.275 ;
      RECT 1303.485 617.545 1303.685 618.275 ;
      RECT 1303.985 617.545 1304.185 618.275 ;
      RECT 1304.48 617.545 1304.68 618.275 ;
      RECT 1304.745 0.3 1305.005 4.63 ;
      RECT 1305.3 617.545 1305.5 618.275 ;
      RECT 1305.765 0.16 1306.535 0.42 ;
      RECT 1305.765 0.16 1306.025 4.63 ;
      RECT 1306.275 0.16 1306.535 8.82 ;
      RECT 1305.255 0.3 1305.515 4.63 ;
      RECT 1305.795 617.545 1305.995 618.275 ;
      RECT 1306.295 617.545 1306.495 618.275 ;
      RECT 1306.795 617.545 1306.995 618.275 ;
      RECT 1307.29 617.545 1307.49 618.275 ;
      RECT 1308.11 617.545 1308.31 618.275 ;
      RECT 1308.605 617.545 1308.805 618.275 ;
      RECT 1309.105 617.545 1309.305 618.275 ;
      RECT 1309.605 617.545 1309.805 618.275 ;
      RECT 1310.1 617.545 1310.3 618.275 ;
      RECT 1310.92 617.545 1311.12 618.275 ;
      RECT 1311.415 617.545 1311.615 618.275 ;
      RECT 1311.915 617.545 1312.115 618.275 ;
      RECT 1312.415 617.545 1312.615 618.275 ;
      RECT 1312.91 617.545 1313.11 618.275 ;
      RECT 1313.73 617.545 1313.93 618.275 ;
      RECT 1314.225 617.545 1314.425 618.275 ;
      RECT 1314.725 617.545 1314.925 618.275 ;
      RECT 1315.225 617.545 1315.425 618.275 ;
      RECT 1315.72 617.545 1315.92 618.275 ;
      RECT 1316.54 617.545 1316.74 618.275 ;
      RECT 1317.035 617.545 1317.235 618.275 ;
      RECT 1317.535 617.545 1317.735 618.275 ;
      RECT 1318.035 617.545 1318.235 618.275 ;
      RECT 1318.53 617.545 1318.73 618.275 ;
      RECT 1319.35 617.545 1319.55 618.275 ;
      RECT 1319.845 617.545 1320.045 618.275 ;
      RECT 1320.045 0.52 1320.305 4.5 ;
      RECT 1320.965 0.165 1321.735 0.425 ;
      RECT 1320.965 0.165 1321.225 8.825 ;
      RECT 1321.475 0.165 1321.735 8.825 ;
      RECT 1320.345 617.545 1320.545 618.275 ;
      RECT 1320.845 617.545 1321.045 618.275 ;
      RECT 1321.34 617.545 1321.54 618.275 ;
      RECT 1321.985 0.3 1322.245 4.63 ;
      RECT 1322.16 617.545 1322.36 618.275 ;
      RECT 1322.495 0.3 1322.755 4.63 ;
      RECT 1322.655 617.545 1322.855 618.275 ;
      RECT 1323.155 617.545 1323.355 618.275 ;
      RECT 1323.655 617.545 1323.855 618.275 ;
      RECT 1324.15 617.545 1324.35 618.275 ;
      RECT 1324.97 617.545 1325.17 618.275 ;
      RECT 1325.465 617.545 1325.665 618.275 ;
      RECT 1325.965 617.545 1326.165 618.275 ;
      RECT 1326.465 617.545 1326.665 618.275 ;
      RECT 1326.96 617.545 1327.16 618.275 ;
      RECT 1327.78 617.545 1327.98 618.275 ;
      RECT 1328.715 0.17 1329.485 0.43 ;
      RECT 1328.715 0.17 1328.975 8.7 ;
      RECT 1329.225 0.17 1329.485 16.7 ;
      RECT 1328.275 617.545 1328.475 618.275 ;
      RECT 1328.775 617.545 1328.975 618.275 ;
      RECT 1329.275 617.545 1329.475 618.275 ;
      RECT 1329.77 617.545 1329.97 618.275 ;
      RECT 1329.735 0.3 1329.995 4.63 ;
      RECT 1330.755 0.17 1331.525 0.43 ;
      RECT 1330.755 0.17 1331.015 8.7 ;
      RECT 1331.265 0.17 1331.525 16.7 ;
      RECT 1330.245 0.3 1330.505 4.63 ;
      RECT 1330.59 617.545 1330.79 618.275 ;
      RECT 1331.085 617.545 1331.285 618.275 ;
      RECT 1331.585 617.545 1331.785 618.275 ;
      RECT 1332.085 617.545 1332.285 618.275 ;
      RECT 1332.58 617.545 1332.78 618.275 ;
      RECT 1333.4 617.545 1333.6 618.275 ;
      RECT 1334.325 0.17 1335.095 0.43 ;
      RECT 1334.325 0.17 1334.585 11.38 ;
      RECT 1334.835 0.17 1335.095 16.7 ;
      RECT 1333.895 617.545 1334.095 618.275 ;
      RECT 1334.395 617.545 1334.595 618.275 ;
      RECT 1334.895 617.545 1335.095 618.275 ;
      RECT 1335.39 617.545 1335.59 618.275 ;
      RECT 1335.7 0.52 1335.96 10.655 ;
      RECT 1336.21 617.545 1336.41 618.275 ;
      RECT 1336.705 617.545 1336.905 618.275 ;
      RECT 1337.205 617.545 1337.405 618.275 ;
      RECT 1337.23 0.52 1337.49 7.94 ;
      RECT 1337.705 617.545 1337.905 618.275 ;
      RECT 1338.2 617.545 1338.4 618.275 ;
      RECT 1339.02 617.545 1339.22 618.275 ;
      RECT 1338.995 0.3 1339.255 8.23 ;
      RECT 1339.515 617.545 1339.715 618.275 ;
      RECT 1340.015 0.165 1340.785 0.425 ;
      RECT 1340.015 0.165 1340.275 8.825 ;
      RECT 1340.525 0.165 1340.785 8.825 ;
      RECT 1339.505 0.3 1339.765 4.63 ;
      RECT 1340.015 617.545 1340.215 618.275 ;
      RECT 1340.515 617.545 1340.715 618.275 ;
      RECT 1341.01 617.545 1341.21 618.275 ;
      RECT 1341.83 617.545 1342.03 618.275 ;
      RECT 1342.325 617.545 1342.525 618.275 ;
      RECT 1342.825 617.545 1343.025 618.275 ;
      RECT 1343.23 0.52 1343.49 4.5 ;
      RECT 1343.325 617.545 1343.525 618.275 ;
      RECT 1343.82 617.545 1344.02 618.275 ;
      RECT 1344.165 0.52 1344.425 10.655 ;
      RECT 1344.64 617.545 1344.84 618.275 ;
      RECT 1345.135 617.545 1345.335 618.275 ;
      RECT 1345.17 0.3 1345.43 4.63 ;
      RECT 1345.635 617.545 1345.835 618.275 ;
      RECT 1346.19 0.16 1346.96 0.42 ;
      RECT 1346.19 0.16 1346.45 8.82 ;
      RECT 1346.7 0.16 1346.96 8.82 ;
      RECT 1345.68 0.3 1345.94 4.63 ;
      RECT 1346.135 617.545 1346.335 618.275 ;
      RECT 1346.63 617.545 1346.83 618.275 ;
      RECT 1347.45 617.545 1347.65 618.275 ;
      RECT 1347.945 617.545 1348.145 618.275 ;
      RECT 1348.445 617.545 1348.645 618.275 ;
      RECT 1348.945 617.545 1349.145 618.275 ;
      RECT 1349.44 617.545 1349.64 618.275 ;
      RECT 1349.705 0.3 1349.965 4.63 ;
      RECT 1350.26 617.545 1350.46 618.275 ;
      RECT 1350.725 0.16 1351.495 0.42 ;
      RECT 1350.725 0.16 1350.985 4.63 ;
      RECT 1351.235 0.16 1351.495 8.82 ;
      RECT 1350.215 0.3 1350.475 4.63 ;
      RECT 1350.755 617.545 1350.955 618.275 ;
      RECT 1351.255 617.545 1351.455 618.275 ;
      RECT 1351.755 617.545 1351.955 618.275 ;
      RECT 1352.25 617.545 1352.45 618.275 ;
      RECT 1353.07 617.545 1353.27 618.275 ;
      RECT 1353.565 617.545 1353.765 618.275 ;
      RECT 1354.065 617.545 1354.265 618.275 ;
      RECT 1354.565 617.545 1354.765 618.275 ;
      RECT 1355.06 617.545 1355.26 618.275 ;
      RECT 1355.88 617.545 1356.08 618.275 ;
      RECT 1356.375 617.545 1356.575 618.275 ;
      RECT 1356.875 617.545 1357.075 618.275 ;
      RECT 1357.375 617.545 1357.575 618.275 ;
      RECT 1357.87 617.545 1358.07 618.275 ;
      RECT 1358.69 617.545 1358.89 618.275 ;
      RECT 1359.185 617.545 1359.385 618.275 ;
      RECT 1359.685 617.545 1359.885 618.275 ;
      RECT 1360.185 617.545 1360.385 618.275 ;
      RECT 1360.68 617.545 1360.88 618.275 ;
      RECT 1361.5 617.545 1361.7 618.275 ;
      RECT 1361.995 617.545 1362.195 618.275 ;
      RECT 1362.495 617.545 1362.695 618.275 ;
      RECT 1362.995 617.545 1363.195 618.275 ;
      RECT 1363.49 617.545 1363.69 618.275 ;
      RECT 1364.31 617.545 1364.51 618.275 ;
      RECT 1364.805 617.545 1365.005 618.275 ;
      RECT 1365.005 0.52 1365.265 4.5 ;
      RECT 1365.925 0.165 1366.695 0.425 ;
      RECT 1365.925 0.165 1366.185 8.825 ;
      RECT 1366.435 0.165 1366.695 8.825 ;
      RECT 1365.305 617.545 1365.505 618.275 ;
      RECT 1365.805 617.545 1366.005 618.275 ;
      RECT 1366.3 617.545 1366.5 618.275 ;
      RECT 1366.945 0.3 1367.205 4.63 ;
      RECT 1367.12 617.545 1367.32 618.275 ;
      RECT 1367.455 0.3 1367.715 4.63 ;
      RECT 1367.615 617.545 1367.815 618.275 ;
      RECT 1368.115 617.545 1368.315 618.275 ;
      RECT 1368.615 617.545 1368.815 618.275 ;
      RECT 1369.11 617.545 1369.31 618.275 ;
      RECT 1369.93 617.545 1370.13 618.275 ;
      RECT 1370.425 617.545 1370.625 618.275 ;
      RECT 1370.925 617.545 1371.125 618.275 ;
      RECT 1371.425 617.545 1371.625 618.275 ;
      RECT 1371.92 617.545 1372.12 618.275 ;
      RECT 1372.74 617.545 1372.94 618.275 ;
      RECT 1373.675 0.17 1374.445 0.43 ;
      RECT 1373.675 0.17 1373.935 8.7 ;
      RECT 1374.185 0.17 1374.445 16.7 ;
      RECT 1373.235 617.545 1373.435 618.275 ;
      RECT 1373.735 617.545 1373.935 618.275 ;
      RECT 1374.235 617.545 1374.435 618.275 ;
      RECT 1374.73 617.545 1374.93 618.275 ;
      RECT 1374.695 0.3 1374.955 4.63 ;
      RECT 1375.715 0.17 1376.485 0.43 ;
      RECT 1375.715 0.17 1375.975 8.7 ;
      RECT 1376.225 0.17 1376.485 16.7 ;
      RECT 1375.205 0.3 1375.465 4.63 ;
      RECT 1375.55 617.545 1375.75 618.275 ;
      RECT 1376.045 617.545 1376.245 618.275 ;
      RECT 1376.545 617.545 1376.745 618.275 ;
      RECT 1377.045 617.545 1377.245 618.275 ;
      RECT 1377.54 617.545 1377.74 618.275 ;
      RECT 1378.36 617.545 1378.56 618.275 ;
      RECT 1379.285 0.17 1380.055 0.43 ;
      RECT 1379.285 0.17 1379.545 11.38 ;
      RECT 1379.795 0.17 1380.055 16.7 ;
      RECT 1378.855 617.545 1379.055 618.275 ;
      RECT 1379.355 617.545 1379.555 618.275 ;
      RECT 1379.855 617.545 1380.055 618.275 ;
      RECT 1380.35 617.545 1380.55 618.275 ;
      RECT 1380.66 0.52 1380.92 10.655 ;
      RECT 1381.17 617.545 1381.37 618.275 ;
      RECT 1381.665 617.545 1381.865 618.275 ;
      RECT 1382.165 617.545 1382.365 618.275 ;
      RECT 1382.19 0.52 1382.45 7.94 ;
      RECT 1382.665 617.545 1382.865 618.275 ;
      RECT 1383.16 617.545 1383.36 618.275 ;
      RECT 1383.98 617.545 1384.18 618.275 ;
      RECT 1383.955 0.3 1384.215 8.23 ;
      RECT 1384.475 617.545 1384.675 618.275 ;
      RECT 1384.975 0.165 1385.745 0.425 ;
      RECT 1384.975 0.165 1385.235 8.825 ;
      RECT 1385.485 0.165 1385.745 8.825 ;
      RECT 1384.465 0.3 1384.725 4.63 ;
      RECT 1384.975 617.545 1385.175 618.275 ;
      RECT 1385.475 617.545 1385.675 618.275 ;
      RECT 1385.97 617.545 1386.17 618.275 ;
      RECT 1386.79 617.545 1386.99 618.275 ;
      RECT 1387.285 617.545 1387.485 618.275 ;
      RECT 1387.785 617.545 1387.985 618.275 ;
      RECT 1388.19 0.52 1388.45 4.5 ;
      RECT 1388.285 617.545 1388.485 618.275 ;
      RECT 1388.78 617.545 1388.98 618.275 ;
      RECT 1389.125 0.52 1389.385 10.655 ;
      RECT 1389.6 617.545 1389.8 618.275 ;
      RECT 1390.095 617.545 1390.295 618.275 ;
      RECT 1390.13 0.3 1390.39 4.63 ;
      RECT 1390.595 617.545 1390.795 618.275 ;
      RECT 1391.15 0.16 1391.92 0.42 ;
      RECT 1391.15 0.16 1391.41 8.82 ;
      RECT 1391.66 0.16 1391.92 8.82 ;
      RECT 1390.64 0.3 1390.9 4.63 ;
      RECT 1391.095 617.545 1391.295 618.275 ;
      RECT 1391.59 617.545 1391.79 618.275 ;
      RECT 1392.41 617.545 1392.61 618.275 ;
      RECT 1392.905 617.545 1393.105 618.275 ;
      RECT 1393.405 617.545 1393.605 618.275 ;
      RECT 1393.905 617.545 1394.105 618.275 ;
      RECT 1394.4 617.545 1394.6 618.275 ;
      RECT 1394.665 0.3 1394.925 4.63 ;
      RECT 1395.22 617.545 1395.42 618.275 ;
      RECT 1395.685 0.16 1396.455 0.42 ;
      RECT 1395.685 0.16 1395.945 4.63 ;
      RECT 1396.195 0.16 1396.455 8.82 ;
      RECT 1395.175 0.3 1395.435 4.63 ;
      RECT 1395.715 617.545 1395.915 618.275 ;
      RECT 1396.215 617.545 1396.415 618.275 ;
      RECT 1396.715 617.545 1396.915 618.275 ;
      RECT 1397.21 617.545 1397.41 618.275 ;
      RECT 1398.03 617.545 1398.23 618.275 ;
      RECT 1398.525 617.545 1398.725 618.275 ;
      RECT 1399.025 617.545 1399.225 618.275 ;
      RECT 1399.525 617.545 1399.725 618.275 ;
      RECT 1400.02 617.545 1400.22 618.275 ;
      RECT 1400.84 617.545 1401.04 618.275 ;
      RECT 1401.335 617.545 1401.535 618.275 ;
      RECT 1401.835 617.545 1402.035 618.275 ;
      RECT 1402.335 617.545 1402.535 618.275 ;
      RECT 1402.83 617.545 1403.03 618.275 ;
      RECT 1403.65 617.545 1403.85 618.275 ;
      RECT 1404.145 617.545 1404.345 618.275 ;
      RECT 1404.645 617.545 1404.845 618.275 ;
      RECT 1405.145 617.545 1405.345 618.275 ;
      RECT 1405.64 617.545 1405.84 618.275 ;
      RECT 1406.46 617.545 1406.66 618.275 ;
      RECT 1406.955 617.545 1407.155 618.275 ;
      RECT 1407.455 617.545 1407.655 618.275 ;
      RECT 1407.955 617.545 1408.155 618.275 ;
      RECT 1408.45 617.545 1408.65 618.275 ;
      RECT 1409.27 617.545 1409.47 618.275 ;
      RECT 1409.765 617.545 1409.965 618.275 ;
      RECT 1409.965 0.52 1410.225 4.5 ;
      RECT 1410.885 0.165 1411.655 0.425 ;
      RECT 1410.885 0.165 1411.145 8.825 ;
      RECT 1411.395 0.165 1411.655 8.825 ;
      RECT 1410.265 617.545 1410.465 618.275 ;
      RECT 1410.765 617.545 1410.965 618.275 ;
      RECT 1411.26 617.545 1411.46 618.275 ;
      RECT 1411.905 0.3 1412.165 4.63 ;
      RECT 1412.08 617.545 1412.28 618.275 ;
      RECT 1412.415 0.3 1412.675 4.63 ;
      RECT 1412.575 617.545 1412.775 618.275 ;
      RECT 1413.075 617.545 1413.275 618.275 ;
      RECT 1413.575 617.545 1413.775 618.275 ;
      RECT 1414.07 617.545 1414.27 618.275 ;
      RECT 1414.89 617.545 1415.09 618.275 ;
      RECT 1415.385 617.545 1415.585 618.275 ;
      RECT 1415.885 617.545 1416.085 618.275 ;
      RECT 1416.385 617.545 1416.585 618.275 ;
      RECT 1416.88 617.545 1417.08 618.275 ;
      RECT 1417.7 617.545 1417.9 618.275 ;
      RECT 1418.635 0.17 1419.405 0.43 ;
      RECT 1418.635 0.17 1418.895 8.7 ;
      RECT 1419.145 0.17 1419.405 16.7 ;
      RECT 1418.195 617.545 1418.395 618.275 ;
      RECT 1418.695 617.545 1418.895 618.275 ;
      RECT 1419.195 617.545 1419.395 618.275 ;
      RECT 1419.69 617.545 1419.89 618.275 ;
      RECT 1419.655 0.3 1419.915 4.63 ;
      RECT 1420.675 0.17 1421.445 0.43 ;
      RECT 1420.675 0.17 1420.935 8.7 ;
      RECT 1421.185 0.17 1421.445 16.7 ;
      RECT 1420.165 0.3 1420.425 4.63 ;
      RECT 1420.51 617.545 1420.71 618.275 ;
      RECT 1421.005 617.545 1421.205 618.275 ;
      RECT 1421.505 617.545 1421.705 618.275 ;
      RECT 1422.005 617.545 1422.205 618.275 ;
      RECT 1422.5 617.545 1422.7 618.275 ;
      RECT 1423.32 617.545 1423.52 618.275 ;
      RECT 1424.245 0.17 1425.015 0.43 ;
      RECT 1424.245 0.17 1424.505 11.38 ;
      RECT 1424.755 0.17 1425.015 16.7 ;
      RECT 1423.815 617.545 1424.015 618.275 ;
      RECT 1424.315 617.545 1424.515 618.275 ;
      RECT 1424.815 617.545 1425.015 618.275 ;
      RECT 1425.31 617.545 1425.51 618.275 ;
      RECT 1425.62 0.52 1425.88 10.655 ;
      RECT 1426.13 617.545 1426.33 618.275 ;
      RECT 1426.625 617.545 1426.825 618.275 ;
      RECT 1427.125 617.545 1427.325 618.275 ;
      RECT 1427.15 0.52 1427.41 7.94 ;
      RECT 1427.625 617.545 1427.825 618.275 ;
      RECT 1428.12 617.545 1428.32 618.275 ;
      RECT 1428.94 617.545 1429.14 618.275 ;
      RECT 1428.915 0.3 1429.175 8.23 ;
      RECT 1429.435 617.545 1429.635 618.275 ;
      RECT 1429.935 0.165 1430.705 0.425 ;
      RECT 1429.935 0.165 1430.195 8.825 ;
      RECT 1430.445 0.165 1430.705 8.825 ;
      RECT 1429.425 0.3 1429.685 4.63 ;
      RECT 1429.935 617.545 1430.135 618.275 ;
      RECT 1430.435 617.545 1430.635 618.275 ;
      RECT 1430.93 617.545 1431.13 618.275 ;
      RECT 1431.75 617.545 1431.95 618.275 ;
      RECT 1432.245 617.545 1432.445 618.275 ;
      RECT 1432.745 617.545 1432.945 618.275 ;
      RECT 1433.15 0.52 1433.41 4.5 ;
      RECT 1433.245 617.545 1433.445 618.275 ;
      RECT 1433.74 617.545 1433.94 618.275 ;
      RECT 1434.085 0.52 1434.345 10.655 ;
      RECT 1434.56 617.545 1434.76 618.275 ;
      RECT 1435.055 617.545 1435.255 618.275 ;
      RECT 1435.09 0.3 1435.35 4.63 ;
      RECT 1435.555 617.545 1435.755 618.275 ;
      RECT 1436.11 0.16 1436.88 0.42 ;
      RECT 1436.11 0.16 1436.37 8.82 ;
      RECT 1436.62 0.16 1436.88 8.82 ;
      RECT 1435.6 0.3 1435.86 4.63 ;
      RECT 1436.055 617.545 1436.255 618.275 ;
      RECT 1436.55 617.545 1436.75 618.275 ;
      RECT 1437.37 617.545 1437.57 618.275 ;
      RECT 1437.865 617.545 1438.065 618.275 ;
      RECT 1438.365 617.545 1438.565 618.275 ;
      RECT 1438.865 617.545 1439.065 618.275 ;
      RECT 1439.36 617.545 1439.56 618.275 ;
      RECT 1439.625 0.3 1439.885 4.63 ;
      RECT 1440.18 617.545 1440.38 618.275 ;
      RECT 1440.645 0.16 1441.415 0.42 ;
      RECT 1440.645 0.16 1440.905 4.63 ;
      RECT 1441.155 0.16 1441.415 8.82 ;
      RECT 1440.135 0.3 1440.395 4.63 ;
      RECT 1440.675 617.545 1440.875 618.275 ;
      RECT 1441.175 617.545 1441.375 618.275 ;
      RECT 1441.675 617.545 1441.875 618.275 ;
      RECT 1442.17 617.545 1442.37 618.275 ;
      RECT 1442.99 617.545 1443.19 618.275 ;
      RECT 1443.485 617.545 1443.685 618.275 ;
      RECT 1443.985 617.545 1444.185 618.275 ;
      RECT 1444.485 617.545 1444.685 618.275 ;
      RECT 1444.98 617.545 1445.18 618.275 ;
      RECT 1445.8 617.545 1446 618.275 ;
      RECT 1446.295 617.545 1446.495 618.275 ;
      RECT 1446.795 617.545 1446.995 618.275 ;
      RECT 1447.295 617.545 1447.495 618.275 ;
      RECT 1447.79 617.545 1447.99 618.275 ;
      RECT 1448.61 617.545 1448.81 618.275 ;
      RECT 1449.105 617.545 1449.305 618.275 ;
      RECT 1449.605 617.545 1449.805 618.275 ;
      RECT 1450.105 617.545 1450.305 618.275 ;
      RECT 1450.6 617.545 1450.8 618.275 ;
      RECT 1451.42 617.545 1451.62 618.275 ;
      RECT 1451.915 617.545 1452.115 618.275 ;
      RECT 1452.415 617.545 1452.615 618.275 ;
      RECT 1452.915 617.545 1453.115 618.275 ;
      RECT 1453.41 617.545 1453.61 618.275 ;
      RECT 1454.23 617.545 1454.43 618.275 ;
      RECT 1454.725 617.545 1454.925 618.275 ;
      RECT 1454.925 0.52 1455.185 4.5 ;
      RECT 1455.845 0.165 1456.615 0.425 ;
      RECT 1455.845 0.165 1456.105 8.825 ;
      RECT 1456.355 0.165 1456.615 8.825 ;
      RECT 1455.225 617.545 1455.425 618.275 ;
      RECT 1455.725 617.545 1455.925 618.275 ;
      RECT 1456.22 617.545 1456.42 618.275 ;
      RECT 1456.865 0.3 1457.125 4.63 ;
      RECT 1457.04 617.545 1457.24 618.275 ;
      RECT 1457.375 0.3 1457.635 4.63 ;
      RECT 1457.535 617.545 1457.735 618.275 ;
      RECT 1458.035 617.545 1458.235 618.275 ;
      RECT 1458.535 617.545 1458.735 618.275 ;
      RECT 1459.03 617.545 1459.23 618.275 ;
      RECT 1459.85 617.545 1460.05 618.275 ;
      RECT 1460.345 617.545 1460.545 618.275 ;
      RECT 1460.845 617.545 1461.045 618.275 ;
      RECT 1461.345 617.545 1461.545 618.275 ;
      RECT 1461.84 617.545 1462.04 618.275 ;
      RECT 1462.66 617.545 1462.86 618.275 ;
      RECT 1463.595 0.17 1464.365 0.43 ;
      RECT 1463.595 0.17 1463.855 8.7 ;
      RECT 1464.105 0.17 1464.365 16.7 ;
      RECT 1463.155 617.545 1463.355 618.275 ;
      RECT 1463.655 617.545 1463.855 618.275 ;
      RECT 1464.155 617.545 1464.355 618.275 ;
      RECT 1464.65 617.545 1464.85 618.275 ;
      RECT 1464.615 0.3 1464.875 4.63 ;
      RECT 1465.635 0.17 1466.405 0.43 ;
      RECT 1465.635 0.17 1465.895 8.7 ;
      RECT 1466.145 0.17 1466.405 16.7 ;
      RECT 1465.125 0.3 1465.385 4.63 ;
      RECT 1465.47 617.545 1465.67 618.275 ;
      RECT 1465.965 617.545 1466.165 618.275 ;
      RECT 1466.465 617.545 1466.665 618.275 ;
      RECT 1466.965 617.545 1467.165 618.275 ;
      RECT 1467.46 617.545 1467.66 618.275 ;
      RECT 1468.28 617.545 1468.48 618.275 ;
      RECT 1469.205 0.17 1469.975 0.43 ;
      RECT 1469.205 0.17 1469.465 11.38 ;
      RECT 1469.715 0.17 1469.975 16.7 ;
      RECT 1468.775 617.545 1468.975 618.275 ;
      RECT 1469.275 617.545 1469.475 618.275 ;
      RECT 1469.775 617.545 1469.975 618.275 ;
      RECT 1470.27 617.545 1470.47 618.275 ;
      RECT 1470.58 0.52 1470.84 10.655 ;
      RECT 1471.09 617.545 1471.29 618.275 ;
      RECT 1471.585 617.545 1471.785 618.275 ;
      RECT 1472.085 617.545 1472.285 618.275 ;
      RECT 1472.11 0.52 1472.37 7.94 ;
      RECT 1472.585 617.545 1472.785 618.275 ;
      RECT 1473.08 617.545 1473.28 618.275 ;
      RECT 1473.9 617.545 1474.1 618.275 ;
      RECT 1473.875 0.3 1474.135 8.23 ;
      RECT 1474.395 617.545 1474.595 618.275 ;
      RECT 1474.895 0.165 1475.665 0.425 ;
      RECT 1474.895 0.165 1475.155 8.825 ;
      RECT 1475.405 0.165 1475.665 8.825 ;
      RECT 1474.385 0.3 1474.645 4.63 ;
      RECT 1474.895 617.545 1475.095 618.275 ;
      RECT 1475.395 617.545 1475.595 618.275 ;
      RECT 1475.89 617.545 1476.09 618.275 ;
      RECT 1476.71 617.545 1476.91 618.275 ;
      RECT 1477.205 617.545 1477.405 618.275 ;
      RECT 1477.705 617.545 1477.905 618.275 ;
      RECT 1478.11 0.52 1478.37 4.5 ;
      RECT 1478.205 617.545 1478.405 618.275 ;
      RECT 1478.7 617.545 1478.9 618.275 ;
      RECT 1479.045 0.52 1479.305 10.655 ;
      RECT 1479.52 617.545 1479.72 618.275 ;
      RECT 1480.015 617.545 1480.215 618.275 ;
      RECT 1480.05 0.3 1480.31 4.63 ;
      RECT 1480.515 617.545 1480.715 618.275 ;
      RECT 1481.07 0.16 1481.84 0.42 ;
      RECT 1481.07 0.16 1481.33 8.82 ;
      RECT 1481.58 0.16 1481.84 8.82 ;
      RECT 1480.56 0.3 1480.82 4.63 ;
      RECT 1481.015 617.545 1481.215 618.275 ;
      RECT 1481.51 617.545 1481.71 618.275 ;
      RECT 1482.33 617.545 1482.53 618.275 ;
      RECT 1482.825 617.545 1483.025 618.275 ;
      RECT 1483.325 617.545 1483.525 618.275 ;
      RECT 1483.825 617.545 1484.025 618.275 ;
      RECT 1484.32 617.545 1484.52 618.275 ;
      RECT 1484.585 0.3 1484.845 4.63 ;
      RECT 1485.14 617.545 1485.34 618.275 ;
      RECT 1485.605 0.16 1486.375 0.42 ;
      RECT 1485.605 0.16 1485.865 4.63 ;
      RECT 1486.115 0.16 1486.375 8.82 ;
      RECT 1485.095 0.3 1485.355 4.63 ;
      RECT 1485.635 617.545 1485.835 618.275 ;
      RECT 1486.135 617.545 1486.335 618.275 ;
      RECT 1486.635 617.545 1486.835 618.275 ;
      RECT 1487.13 617.545 1487.33 618.275 ;
      RECT 1487.95 617.545 1488.15 618.275 ;
      RECT 1488.445 617.545 1488.645 618.275 ;
      RECT 1488.945 617.545 1489.145 618.275 ;
      RECT 1489.445 617.545 1489.645 618.275 ;
      RECT 1489.94 617.545 1490.14 618.275 ;
      RECT 1490.76 617.545 1490.96 618.275 ;
      RECT 1491.255 617.545 1491.455 618.275 ;
      RECT 1491.755 617.545 1491.955 618.275 ;
      RECT 1492.255 617.545 1492.455 618.275 ;
      RECT 1492.75 617.545 1492.95 618.275 ;
      RECT 1493.57 617.545 1493.77 618.275 ;
      RECT 1494.065 617.545 1494.265 618.275 ;
      RECT 1494.565 617.545 1494.765 618.275 ;
      RECT 1495.065 617.545 1495.265 618.275 ;
      RECT 1495.56 617.545 1495.76 618.275 ;
      RECT 1496.38 617.545 1496.58 618.275 ;
      RECT 1496.875 617.545 1497.075 618.275 ;
      RECT 1497.375 617.545 1497.575 618.275 ;
      RECT 1497.875 617.545 1498.075 618.275 ;
      RECT 1498.37 617.545 1498.57 618.275 ;
      RECT 1499.19 617.545 1499.39 618.275 ;
      RECT 1499.685 617.545 1499.885 618.275 ;
      RECT 1499.885 0.52 1500.145 4.5 ;
      RECT 1500.805 0.165 1501.575 0.425 ;
      RECT 1500.805 0.165 1501.065 8.825 ;
      RECT 1501.315 0.165 1501.575 8.825 ;
      RECT 1500.185 617.545 1500.385 618.275 ;
      RECT 1500.685 617.545 1500.885 618.275 ;
      RECT 1501.18 617.545 1501.38 618.275 ;
      RECT 1501.825 0.3 1502.085 4.63 ;
      RECT 1502 617.545 1502.2 618.275 ;
      RECT 1502.335 0.3 1502.595 4.63 ;
      RECT 1502.495 617.545 1502.695 618.275 ;
      RECT 1502.995 617.545 1503.195 618.275 ;
      RECT 1503.495 617.545 1503.695 618.275 ;
      RECT 1503.99 617.545 1504.19 618.275 ;
      RECT 1504.81 617.545 1505.01 618.275 ;
      RECT 1505.305 617.545 1505.505 618.275 ;
      RECT 1505.805 617.545 1506.005 618.275 ;
      RECT 1506.305 617.545 1506.505 618.275 ;
      RECT 1506.8 617.545 1507 618.275 ;
      RECT 1507.62 617.545 1507.82 618.275 ;
      RECT 1508.555 0.17 1509.325 0.43 ;
      RECT 1508.555 0.17 1508.815 8.7 ;
      RECT 1509.065 0.17 1509.325 16.7 ;
      RECT 1508.115 617.545 1508.315 618.275 ;
      RECT 1508.615 617.545 1508.815 618.275 ;
      RECT 1509.115 617.545 1509.315 618.275 ;
      RECT 1509.61 617.545 1509.81 618.275 ;
      RECT 1509.575 0.3 1509.835 4.63 ;
      RECT 1510.595 0.17 1511.365 0.43 ;
      RECT 1510.595 0.17 1510.855 8.7 ;
      RECT 1511.105 0.17 1511.365 16.7 ;
      RECT 1510.085 0.3 1510.345 4.63 ;
      RECT 1510.43 617.545 1510.63 618.275 ;
      RECT 1510.925 617.545 1511.125 618.275 ;
      RECT 1511.425 617.545 1511.625 618.275 ;
      RECT 1511.925 617.545 1512.125 618.275 ;
      RECT 1512.42 617.545 1512.62 618.275 ;
      RECT 1513.24 617.545 1513.44 618.275 ;
      RECT 1514.165 0.17 1514.935 0.43 ;
      RECT 1514.165 0.17 1514.425 11.38 ;
      RECT 1514.675 0.17 1514.935 16.7 ;
      RECT 1513.735 617.545 1513.935 618.275 ;
      RECT 1514.235 617.545 1514.435 618.275 ;
      RECT 1514.735 617.545 1514.935 618.275 ;
      RECT 1515.23 617.545 1515.43 618.275 ;
      RECT 1515.54 0.52 1515.8 10.655 ;
      RECT 1516.05 617.545 1516.25 618.275 ;
      RECT 1516.545 617.545 1516.745 618.275 ;
      RECT 1517.045 617.545 1517.245 618.275 ;
      RECT 1517.07 0.52 1517.33 7.94 ;
      RECT 1517.545 617.545 1517.745 618.275 ;
      RECT 1518.04 617.545 1518.24 618.275 ;
      RECT 1518.86 617.545 1519.06 618.275 ;
      RECT 1519.855 37.065 1520.055 618.275 ;
    LAYER Metal2 SPACING 0.21 ;
      RECT 632.79 0 633.54 618.3 ;
      RECT 626.79 0 632.01 618.3 ;
      RECT 605.015 0 625.075 618.3 ;
      RECT 589.36 0 604.235 618.3 ;
      RECT 587.83 0 588.58 618.3 ;
      RECT 581.83 0 587.05 618.3 ;
      RECT 560.055 0 580.115 618.3 ;
      RECT 544.4 0 559.275 618.3 ;
      RECT 542.87 0 543.62 618.3 ;
      RECT 536.87 0 542.09 618.3 ;
      RECT 515.095 0 535.155 618.3 ;
      RECT 499.44 0 514.315 618.3 ;
      RECT 497.91 0 498.66 618.3 ;
      RECT 491.91 0 497.13 618.3 ;
      RECT 470.135 0 490.195 618.3 ;
      RECT 454.48 0 469.355 618.3 ;
      RECT 452.95 0 453.7 618.3 ;
      RECT 446.95 0 452.17 618.3 ;
      RECT 425.175 0 445.235 618.3 ;
      RECT 409.52 0 424.395 618.3 ;
      RECT 407.99 0 408.74 618.3 ;
      RECT 401.99 0 407.21 618.3 ;
      RECT 380.215 0 400.275 618.3 ;
      RECT 364.56 0 379.435 618.3 ;
      RECT 363.03 0 363.78 618.3 ;
      RECT 357.03 0 362.25 618.3 ;
      RECT 335.255 0 355.315 618.3 ;
      RECT 319.6 0 334.475 618.3 ;
      RECT 318.07 0 318.82 618.3 ;
      RECT 312.07 0 317.29 618.3 ;
      RECT 290.295 0 310.355 618.3 ;
      RECT 274.64 0 289.515 618.3 ;
      RECT 273.11 0 273.86 618.3 ;
      RECT 267.11 0 272.33 618.3 ;
      RECT 245.335 0 265.395 618.3 ;
      RECT 229.68 0 244.555 618.3 ;
      RECT 228.15 0 228.9 618.3 ;
      RECT 222.15 0 227.37 618.3 ;
      RECT 200.375 0 220.435 618.3 ;
      RECT 184.72 0 199.595 618.3 ;
      RECT 183.19 0 183.94 618.3 ;
      RECT 177.19 0 182.41 618.3 ;
      RECT 155.415 0 175.475 618.3 ;
      RECT 139.76 0 154.635 618.3 ;
      RECT 138.23 0 138.98 618.3 ;
      RECT 132.23 0 137.45 618.3 ;
      RECT 110.455 0 130.515 618.3 ;
      RECT 94.8 0 109.675 618.3 ;
      RECT 93.27 0 94.02 618.3 ;
      RECT 87.27 0 92.49 618.3 ;
      RECT 65.495 0 85.555 618.3 ;
      RECT 49.84 0 64.715 618.3 ;
      RECT 48.31 0 49.06 618.3 ;
      RECT 42.31 0 47.53 618.3 ;
      RECT 20.535 0 40.595 618.3 ;
      RECT 4.88 0 19.755 618.3 ;
      RECT 3.35 0 4.1 618.3 ;
      RECT 0 0 2.57 618.3 ;
      RECT 0 0.52 1520.16 618.3 ;
      RECT 1517.59 0 1520.16 618.3 ;
      RECT 1516.06 0 1516.81 618.3 ;
      RECT 1500.405 0 1515.28 618.3 ;
      RECT 1479.565 0 1499.625 618.3 ;
      RECT 1472.63 0 1477.85 618.3 ;
      RECT 1471.1 0 1471.85 618.3 ;
      RECT 1455.445 0 1470.32 618.3 ;
      RECT 1434.605 0 1454.665 618.3 ;
      RECT 1427.67 0 1432.89 618.3 ;
      RECT 1426.14 0 1426.89 618.3 ;
      RECT 1410.485 0 1425.36 618.3 ;
      RECT 1389.645 0 1409.705 618.3 ;
      RECT 1382.71 0 1387.93 618.3 ;
      RECT 1381.18 0 1381.93 618.3 ;
      RECT 1365.525 0 1380.4 618.3 ;
      RECT 1344.685 0 1364.745 618.3 ;
      RECT 1337.75 0 1342.97 618.3 ;
      RECT 1336.22 0 1336.97 618.3 ;
      RECT 1320.565 0 1335.44 618.3 ;
      RECT 1299.725 0 1319.785 618.3 ;
      RECT 1292.79 0 1298.01 618.3 ;
      RECT 1291.26 0 1292.01 618.3 ;
      RECT 1275.605 0 1290.48 618.3 ;
      RECT 1254.765 0 1274.825 618.3 ;
      RECT 1247.83 0 1253.05 618.3 ;
      RECT 1246.3 0 1247.05 618.3 ;
      RECT 1230.645 0 1245.52 618.3 ;
      RECT 1209.805 0 1229.865 618.3 ;
      RECT 1202.87 0 1208.09 618.3 ;
      RECT 1201.34 0 1202.09 618.3 ;
      RECT 1185.685 0 1200.56 618.3 ;
      RECT 1164.845 0 1184.905 618.3 ;
      RECT 1157.91 0 1163.13 618.3 ;
      RECT 1156.38 0 1157.13 618.3 ;
      RECT 1140.725 0 1155.6 618.3 ;
      RECT 1119.885 0 1139.945 618.3 ;
      RECT 1112.95 0 1118.17 618.3 ;
      RECT 1111.42 0 1112.17 618.3 ;
      RECT 1095.765 0 1110.64 618.3 ;
      RECT 1074.925 0 1094.985 618.3 ;
      RECT 1067.99 0 1073.21 618.3 ;
      RECT 1066.46 0 1067.21 618.3 ;
      RECT 1050.805 0 1065.68 618.3 ;
      RECT 1029.965 0 1050.025 618.3 ;
      RECT 1023.03 0 1028.25 618.3 ;
      RECT 1021.5 0 1022.25 618.3 ;
      RECT 1005.845 0 1020.72 618.3 ;
      RECT 985.005 0 1005.065 618.3 ;
      RECT 978.07 0 983.29 618.3 ;
      RECT 976.54 0 977.29 618.3 ;
      RECT 960.885 0 975.76 618.3 ;
      RECT 940.045 0 960.105 618.3 ;
      RECT 933.11 0 938.33 618.3 ;
      RECT 931.58 0 932.33 618.3 ;
      RECT 915.925 0 930.8 618.3 ;
      RECT 895.085 0 915.145 618.3 ;
      RECT 888.15 0 893.37 618.3 ;
      RECT 886.62 0 887.37 618.3 ;
      RECT 870.965 0 885.84 618.3 ;
      RECT 850.125 0 870.185 618.3 ;
      RECT 843.19 0 848.41 618.3 ;
      RECT 841.66 0 842.41 618.3 ;
      RECT 826.005 0 840.88 618.3 ;
      RECT 805.165 0 825.225 618.3 ;
      RECT 776.68 0.17 803.45 618.3 ;
      RECT 776.69 0 803.45 618.3 ;
      RECT 775.16 0 775.91 618.3 ;
      RECT 770.06 0 773.87 618.3 ;
      RECT 768.02 0 768.77 618.3 ;
      RECT 761.39 0 762.65 618.3 ;
      RECT 759.86 0 760.1 618.3 ;
      RECT 758.33 0 758.57 618.3 ;
      RECT 755.27 0 755.51 618.3 ;
      RECT 753.74 0 753.98 618.3 ;
      RECT 747.11 0 752.45 618.3 ;
      RECT 743.53 0 743.79 618.3 ;
      RECT 742.01 0 742.76 618.3 ;
      RECT 716.71 0 741.24 618.3 ;
      RECT 694.935 0 714.995 618.3 ;
      RECT 679.28 0 694.155 618.3 ;
      RECT 677.75 0 678.5 618.3 ;
      RECT 671.75 0 676.97 618.3 ;
      RECT 649.975 0 670.035 618.3 ;
      RECT 634.32 0 649.195 618.3 ;
    LAYER Metal3 ;
      RECT 0 0 1520.16 618.3 ;
    LAYER Metal4 ;
      RECT 4.26 599.405 7.07 618.3 ;
      RECT 4.26 0 7.07 30.425 ;
      RECT 9.88 599.405 12.69 618.3 ;
      RECT 9.88 0 12.69 37.065 ;
      RECT 49.22 599.405 52.03 618.3 ;
      RECT 49.22 0 52.03 30.425 ;
      RECT 54.84 599.405 57.65 618.3 ;
      RECT 54.84 0 57.65 37.065 ;
      RECT 94.18 599.405 96.99 618.3 ;
      RECT 94.18 0 96.99 30.425 ;
      RECT 99.8 599.405 102.61 618.3 ;
      RECT 99.8 0 102.61 37.065 ;
      RECT 139.14 599.405 141.95 618.3 ;
      RECT 139.14 0 141.95 30.425 ;
      RECT 144.76 599.405 147.57 618.3 ;
      RECT 144.76 0 147.57 37.065 ;
      RECT 184.1 599.405 186.91 618.3 ;
      RECT 184.1 0 186.91 30.425 ;
      RECT 189.72 599.405 192.53 618.3 ;
      RECT 189.72 0 192.53 37.065 ;
      RECT 229.06 599.405 231.87 618.3 ;
      RECT 229.06 0 231.87 30.425 ;
      RECT 234.68 599.405 237.49 618.3 ;
      RECT 234.68 0 237.49 37.065 ;
      RECT 274.02 599.405 276.83 618.3 ;
      RECT 274.02 0 276.83 30.425 ;
      RECT 279.64 599.405 282.45 618.3 ;
      RECT 279.64 0 282.45 37.065 ;
      RECT 318.98 599.405 321.79 618.3 ;
      RECT 318.98 0 321.79 30.425 ;
      RECT 324.6 599.405 327.41 618.3 ;
      RECT 324.6 0 327.41 37.065 ;
      RECT 363.94 599.405 366.75 618.3 ;
      RECT 363.94 0 366.75 30.425 ;
      RECT 369.56 599.405 372.37 618.3 ;
      RECT 369.56 0 372.37 37.065 ;
      RECT 408.9 599.405 411.71 618.3 ;
      RECT 408.9 0 411.71 30.425 ;
      RECT 414.52 599.405 417.33 618.3 ;
      RECT 414.52 0 417.33 37.065 ;
      RECT 453.86 599.405 456.67 618.3 ;
      RECT 453.86 0 456.67 30.425 ;
      RECT 459.48 599.405 462.29 618.3 ;
      RECT 459.48 0 462.29 37.065 ;
      RECT 498.82 599.405 501.63 618.3 ;
      RECT 498.82 0 501.63 30.425 ;
      RECT 504.44 599.405 507.25 618.3 ;
      RECT 504.44 0 507.25 37.065 ;
      RECT 543.78 599.405 546.59 618.3 ;
      RECT 543.78 0 546.59 30.425 ;
      RECT 549.4 599.405 552.21 618.3 ;
      RECT 549.4 0 552.21 37.065 ;
      RECT 588.74 599.405 591.55 618.3 ;
      RECT 588.74 0 591.55 30.425 ;
      RECT 594.36 599.405 597.17 618.3 ;
      RECT 594.36 0 597.17 37.065 ;
      RECT 633.7 599.405 636.51 618.3 ;
      RECT 633.7 0 636.51 30.425 ;
      RECT 639.32 599.405 642.13 618.3 ;
      RECT 639.32 0 642.13 37.065 ;
      RECT 678.66 599.405 681.47 618.3 ;
      RECT 678.66 0 681.47 30.425 ;
      RECT 684.28 599.405 687.09 618.3 ;
      RECT 684.28 0 687.09 37.065 ;
      RECT 833.07 599.405 835.88 618.3 ;
      RECT 833.07 0 835.88 37.065 ;
      RECT 838.69 599.405 841.5 618.3 ;
    LAYER Metal4 SPACING 0.21 ;
      RECT 779.77 0 799.09 618.3 ;
      RECT 774.62 0 776.44 618.3 ;
      RECT 769.47 0 771.29 618.3 ;
      RECT 1504.92 0 1520.16 618.3 ;
      RECT 1499.3 0 1501.59 618.3 ;
      RECT 1499.3 30.685 1520.16 36.805 ;
      RECT 1493.68 0 1495.97 618.3 ;
      RECT 1488.06 0 1490.35 618.3 ;
      RECT 1488.06 30.685 1495.97 36.805 ;
      RECT 1482.44 0 1484.73 618.3 ;
      RECT 1476.82 0 1479.11 618.3 ;
      RECT 1476.82 30.685 1484.73 36.805 ;
      RECT 1459.96 0 1473.49 618.3 ;
      RECT 1454.34 0 1456.63 618.3 ;
      RECT 1454.34 30.685 1473.49 36.805 ;
      RECT 1448.72 0 1451.01 618.3 ;
      RECT 1443.1 0 1445.39 618.3 ;
      RECT 1443.1 30.685 1451.01 36.805 ;
      RECT 1437.48 0 1439.77 618.3 ;
      RECT 1431.86 0 1434.15 618.3 ;
      RECT 1431.86 30.685 1439.77 36.805 ;
      RECT 1415 0 1428.53 618.3 ;
      RECT 1409.38 0 1411.67 618.3 ;
      RECT 1409.38 30.685 1428.53 36.805 ;
      RECT 1403.76 0 1406.05 618.3 ;
      RECT 1398.14 0 1400.43 618.3 ;
      RECT 1398.14 30.685 1406.05 36.805 ;
      RECT 1392.52 0 1394.81 618.3 ;
      RECT 1386.9 0 1389.19 618.3 ;
      RECT 1386.9 30.685 1394.81 36.805 ;
      RECT 1370.04 0 1383.57 618.3 ;
      RECT 1364.42 0 1366.71 618.3 ;
      RECT 1364.42 30.685 1383.57 36.805 ;
      RECT 1358.8 0 1361.09 618.3 ;
      RECT 1353.18 0 1355.47 618.3 ;
      RECT 1353.18 30.685 1361.09 36.805 ;
      RECT 1347.56 0 1349.85 618.3 ;
      RECT 1341.94 0 1344.23 618.3 ;
      RECT 1341.94 30.685 1349.85 36.805 ;
      RECT 1325.08 0 1338.61 618.3 ;
      RECT 1319.46 0 1321.75 618.3 ;
      RECT 1319.46 30.685 1338.61 36.805 ;
      RECT 1313.84 0 1316.13 618.3 ;
      RECT 1308.22 0 1310.51 618.3 ;
      RECT 1308.22 30.685 1316.13 36.805 ;
      RECT 1302.6 0 1304.89 618.3 ;
      RECT 1296.98 0 1299.27 618.3 ;
      RECT 1296.98 30.685 1304.89 36.805 ;
      RECT 1280.12 0 1293.65 618.3 ;
      RECT 1274.5 0 1276.79 618.3 ;
      RECT 1274.5 30.685 1293.65 36.805 ;
      RECT 1268.88 0 1271.17 618.3 ;
      RECT 1263.26 0 1265.55 618.3 ;
      RECT 1263.26 30.685 1271.17 36.805 ;
      RECT 1257.64 0 1259.93 618.3 ;
      RECT 1252.02 0 1254.31 618.3 ;
      RECT 1252.02 30.685 1259.93 36.805 ;
      RECT 1235.16 0 1248.69 618.3 ;
      RECT 1229.54 0 1231.83 618.3 ;
      RECT 1229.54 30.685 1248.69 36.805 ;
      RECT 1223.92 0 1226.21 618.3 ;
      RECT 1218.3 0 1220.59 618.3 ;
      RECT 1218.3 30.685 1226.21 36.805 ;
      RECT 1212.68 0 1214.97 618.3 ;
      RECT 1207.06 0 1209.35 618.3 ;
      RECT 1207.06 30.685 1214.97 36.805 ;
      RECT 614.29 0 616.58 618.3 ;
      RECT 608.67 0 610.96 618.3 ;
      RECT 608.67 30.685 616.58 36.805 ;
      RECT 603.05 0 605.34 618.3 ;
      RECT 586.19 0 599.72 618.3 ;
      RECT 586.19 30.685 605.34 36.805 ;
      RECT 580.57 0 582.86 618.3 ;
      RECT 574.95 0 577.24 618.3 ;
      RECT 574.95 30.685 582.86 36.805 ;
      RECT 569.33 0 571.62 618.3 ;
      RECT 563.71 0 566 618.3 ;
      RECT 563.71 30.685 571.62 36.805 ;
      RECT 558.09 0 560.38 618.3 ;
      RECT 541.23 0 554.76 618.3 ;
      RECT 541.23 30.685 560.38 36.805 ;
      RECT 535.61 0 537.9 618.3 ;
      RECT 529.99 0 532.28 618.3 ;
      RECT 529.99 30.685 537.9 36.805 ;
      RECT 524.37 0 526.66 618.3 ;
      RECT 518.75 0 521.04 618.3 ;
      RECT 518.75 30.685 526.66 36.805 ;
      RECT 513.13 0 515.42 618.3 ;
      RECT 496.27 0 509.8 618.3 ;
      RECT 496.27 30.685 515.42 36.805 ;
      RECT 490.65 0 492.94 618.3 ;
      RECT 485.03 0 487.32 618.3 ;
      RECT 485.03 30.685 492.94 36.805 ;
      RECT 479.41 0 481.7 618.3 ;
      RECT 473.79 0 476.08 618.3 ;
      RECT 473.79 30.685 481.7 36.805 ;
      RECT 468.17 0 470.46 618.3 ;
      RECT 451.31 0 464.84 618.3 ;
      RECT 451.31 30.685 470.46 36.805 ;
      RECT 445.69 0 447.98 618.3 ;
      RECT 440.07 0 442.36 618.3 ;
      RECT 440.07 30.685 447.98 36.805 ;
      RECT 434.45 0 436.74 618.3 ;
      RECT 428.83 0 431.12 618.3 ;
      RECT 428.83 30.685 436.74 36.805 ;
      RECT 423.21 0 425.5 618.3 ;
      RECT 406.35 0 419.88 618.3 ;
      RECT 406.35 30.685 425.5 36.805 ;
      RECT 400.73 0 403.02 618.3 ;
      RECT 395.11 0 397.4 618.3 ;
      RECT 395.11 30.685 403.02 36.805 ;
      RECT 389.49 0 391.78 618.3 ;
      RECT 383.87 0 386.16 618.3 ;
      RECT 383.87 30.685 391.78 36.805 ;
      RECT 378.25 0 380.54 618.3 ;
      RECT 361.39 0 374.92 618.3 ;
      RECT 361.39 30.685 380.54 36.805 ;
      RECT 355.77 0 358.06 618.3 ;
      RECT 350.15 0 352.44 618.3 ;
      RECT 350.15 30.685 358.06 36.805 ;
      RECT 344.53 0 346.82 618.3 ;
      RECT 338.91 0 341.2 618.3 ;
      RECT 338.91 30.685 346.82 36.805 ;
      RECT 333.29 0 335.58 618.3 ;
      RECT 316.43 0 329.96 618.3 ;
      RECT 316.43 30.685 335.58 36.805 ;
      RECT 310.81 0 313.1 618.3 ;
      RECT 305.19 0 307.48 618.3 ;
      RECT 305.19 30.685 313.1 36.805 ;
      RECT 299.57 0 301.86 618.3 ;
      RECT 293.95 0 296.24 618.3 ;
      RECT 293.95 30.685 301.86 36.805 ;
      RECT 288.33 0 290.62 618.3 ;
      RECT 271.47 0 285 618.3 ;
      RECT 271.47 30.685 290.62 36.805 ;
      RECT 265.85 0 268.14 618.3 ;
      RECT 260.23 0 262.52 618.3 ;
      RECT 260.23 30.685 268.14 36.805 ;
      RECT 254.61 0 256.9 618.3 ;
      RECT 248.99 0 251.28 618.3 ;
      RECT 248.99 30.685 256.9 36.805 ;
      RECT 243.37 0 245.66 618.3 ;
      RECT 226.51 0 240.04 618.3 ;
      RECT 226.51 30.685 245.66 36.805 ;
      RECT 220.89 0 223.18 618.3 ;
      RECT 215.27 0 217.56 618.3 ;
      RECT 215.27 30.685 223.18 36.805 ;
      RECT 209.65 0 211.94 618.3 ;
      RECT 204.03 0 206.32 618.3 ;
      RECT 204.03 30.685 211.94 36.805 ;
      RECT 198.41 0 200.7 618.3 ;
      RECT 181.55 0 195.08 618.3 ;
      RECT 181.55 30.685 200.7 36.805 ;
      RECT 175.93 0 178.22 618.3 ;
      RECT 170.31 0 172.6 618.3 ;
      RECT 170.31 30.685 178.22 36.805 ;
      RECT 164.69 0 166.98 618.3 ;
      RECT 159.07 0 161.36 618.3 ;
      RECT 159.07 30.685 166.98 36.805 ;
      RECT 153.45 0 155.74 618.3 ;
      RECT 136.59 0 150.12 618.3 ;
      RECT 136.59 30.685 155.74 36.805 ;
      RECT 130.97 0 133.26 618.3 ;
      RECT 125.35 0 127.64 618.3 ;
      RECT 125.35 30.685 133.26 36.805 ;
      RECT 119.73 0 122.02 618.3 ;
      RECT 114.11 0 116.4 618.3 ;
      RECT 114.11 30.685 122.02 36.805 ;
      RECT 108.49 0 110.78 618.3 ;
      RECT 91.63 0 105.16 618.3 ;
      RECT 91.63 30.685 110.78 36.805 ;
      RECT 86.01 0 88.3 618.3 ;
      RECT 80.39 0 82.68 618.3 ;
      RECT 80.39 30.685 88.3 36.805 ;
      RECT 74.77 0 77.06 618.3 ;
      RECT 69.15 0 71.44 618.3 ;
      RECT 69.15 30.685 77.06 36.805 ;
      RECT 63.53 0 65.82 618.3 ;
      RECT 46.67 0 60.2 618.3 ;
      RECT 46.67 30.685 65.82 36.805 ;
      RECT 41.05 0 43.34 618.3 ;
      RECT 35.43 0 37.72 618.3 ;
      RECT 35.43 30.685 43.34 36.805 ;
      RECT 29.81 0 32.1 618.3 ;
      RECT 24.19 0 26.48 618.3 ;
      RECT 24.19 30.685 32.1 36.805 ;
      RECT 18.57 0 20.86 618.3 ;
      RECT 0 0 15.24 618.3 ;
      RECT 0 30.685 20.86 36.805 ;
      RECT 1190.2 0 1203.73 618.3 ;
      RECT 1184.58 0 1186.87 618.3 ;
      RECT 1184.58 30.685 1203.73 36.805 ;
      RECT 1178.96 0 1181.25 618.3 ;
      RECT 1173.34 0 1175.63 618.3 ;
      RECT 1173.34 30.685 1181.25 36.805 ;
      RECT 1167.72 0 1170.01 618.3 ;
      RECT 1162.1 0 1164.39 618.3 ;
      RECT 1162.1 30.685 1170.01 36.805 ;
      RECT 1145.24 0 1158.77 618.3 ;
      RECT 1139.62 0 1141.91 618.3 ;
      RECT 1139.62 30.685 1158.77 36.805 ;
      RECT 1134 0 1136.29 618.3 ;
      RECT 1128.38 0 1130.67 618.3 ;
      RECT 1128.38 30.685 1136.29 36.805 ;
      RECT 1122.76 0 1125.05 618.3 ;
      RECT 1117.14 0 1119.43 618.3 ;
      RECT 1117.14 30.685 1125.05 36.805 ;
      RECT 1100.28 0 1113.81 618.3 ;
      RECT 1094.66 0 1096.95 618.3 ;
      RECT 1094.66 30.685 1113.81 36.805 ;
      RECT 1089.04 0 1091.33 618.3 ;
      RECT 1083.42 0 1085.71 618.3 ;
      RECT 1083.42 30.685 1091.33 36.805 ;
      RECT 1077.8 0 1080.09 618.3 ;
      RECT 1072.18 0 1074.47 618.3 ;
      RECT 1072.18 30.685 1080.09 36.805 ;
      RECT 1055.32 0 1068.85 618.3 ;
      RECT 1049.7 0 1051.99 618.3 ;
      RECT 1049.7 30.685 1068.85 36.805 ;
      RECT 1044.08 0 1046.37 618.3 ;
      RECT 1038.46 0 1040.75 618.3 ;
      RECT 1038.46 30.685 1046.37 36.805 ;
      RECT 1032.84 0 1035.13 618.3 ;
      RECT 1027.22 0 1029.51 618.3 ;
      RECT 1027.22 30.685 1035.13 36.805 ;
      RECT 1010.36 0 1023.89 618.3 ;
      RECT 1004.74 0 1007.03 618.3 ;
      RECT 1004.74 30.685 1023.89 36.805 ;
      RECT 999.12 0 1001.41 618.3 ;
      RECT 993.5 0 995.79 618.3 ;
      RECT 993.5 30.685 1001.41 36.805 ;
      RECT 987.88 0 990.17 618.3 ;
      RECT 982.26 0 984.55 618.3 ;
      RECT 982.26 30.685 990.17 36.805 ;
      RECT 965.4 0 978.93 618.3 ;
      RECT 959.78 0 962.07 618.3 ;
      RECT 959.78 30.685 978.93 36.805 ;
      RECT 954.16 0 956.45 618.3 ;
      RECT 948.54 0 950.83 618.3 ;
      RECT 948.54 30.685 956.45 36.805 ;
      RECT 942.92 0 945.21 618.3 ;
      RECT 937.3 0 939.59 618.3 ;
      RECT 937.3 30.685 945.21 36.805 ;
      RECT 920.44 0 933.97 618.3 ;
      RECT 914.82 0 917.11 618.3 ;
      RECT 914.82 30.685 933.97 36.805 ;
      RECT 909.2 0 911.49 618.3 ;
      RECT 903.58 0 905.87 618.3 ;
      RECT 903.58 30.685 911.49 36.805 ;
      RECT 897.96 0 900.25 618.3 ;
      RECT 892.34 0 894.63 618.3 ;
      RECT 892.34 30.685 900.25 36.805 ;
      RECT 875.48 0 889.01 618.3 ;
      RECT 869.86 0 872.15 618.3 ;
      RECT 869.86 30.685 889.01 36.805 ;
      RECT 864.24 0 866.53 618.3 ;
      RECT 858.62 0 860.91 618.3 ;
      RECT 858.62 30.685 866.53 36.805 ;
      RECT 853 0 855.29 618.3 ;
      RECT 847.38 0 849.67 618.3 ;
      RECT 847.38 30.685 855.29 36.805 ;
      RECT 830.52 0 844.05 618.3 ;
      RECT 824.9 0 827.19 618.3 ;
      RECT 824.9 30.685 844.05 36.805 ;
      RECT 819.28 0 821.57 618.3 ;
      RECT 813.66 0 815.95 618.3 ;
      RECT 813.66 30.685 821.57 36.805 ;
      RECT 808.04 0 810.33 618.3 ;
      RECT 802.42 0 804.71 618.3 ;
      RECT 802.42 30.685 810.33 36.805 ;
      RECT 764.32 0 766.14 618.3 ;
      RECT 759.17 0 760.99 618.3 ;
      RECT 754.02 0 755.84 618.3 ;
      RECT 748.87 0 750.69 618.3 ;
      RECT 743.72 0 745.54 618.3 ;
      RECT 721.07 0 740.39 618.3 ;
      RECT 715.45 0 717.74 618.3 ;
      RECT 709.83 0 712.12 618.3 ;
      RECT 709.83 30.685 717.74 36.805 ;
      RECT 704.21 0 706.5 618.3 ;
      RECT 698.59 0 700.88 618.3 ;
      RECT 698.59 30.685 706.5 36.805 ;
      RECT 692.97 0 695.26 618.3 ;
      RECT 676.11 0 689.64 618.3 ;
      RECT 676.11 30.685 695.26 36.805 ;
      RECT 670.49 0 672.78 618.3 ;
      RECT 664.87 0 667.16 618.3 ;
      RECT 664.87 30.685 672.78 36.805 ;
      RECT 659.25 0 661.54 618.3 ;
      RECT 653.63 0 655.92 618.3 ;
      RECT 653.63 30.685 661.54 36.805 ;
      RECT 648.01 0 650.3 618.3 ;
      RECT 631.15 0 644.68 618.3 ;
      RECT 631.15 30.685 650.3 36.805 ;
      RECT 625.53 0 627.82 618.3 ;
      RECT 619.91 0 622.2 618.3 ;
      RECT 619.91 30.685 627.82 36.805 ;
    LAYER Metal4 ;
      RECT 1513.09 0 1515.9 30.425 ;
      RECT 1513.09 599.405 1515.9 618.3 ;
      RECT 1507.47 0 1510.28 37.065 ;
      RECT 1507.47 599.405 1510.28 618.3 ;
      RECT 1468.13 0 1470.94 30.425 ;
      RECT 1468.13 599.405 1470.94 618.3 ;
      RECT 1462.51 0 1465.32 37.065 ;
      RECT 1462.51 599.405 1465.32 618.3 ;
      RECT 1423.17 0 1425.98 30.425 ;
      RECT 1423.17 599.405 1425.98 618.3 ;
      RECT 1417.55 0 1420.36 37.065 ;
      RECT 1417.55 599.405 1420.36 618.3 ;
      RECT 1378.21 0 1381.02 30.425 ;
      RECT 1378.21 599.405 1381.02 618.3 ;
      RECT 1372.59 0 1375.4 37.065 ;
      RECT 1372.59 599.405 1375.4 618.3 ;
      RECT 1333.25 0 1336.06 30.425 ;
      RECT 1333.25 599.405 1336.06 618.3 ;
      RECT 1327.63 0 1330.44 37.065 ;
      RECT 1327.63 599.405 1330.44 618.3 ;
      RECT 1288.29 0 1291.1 30.425 ;
      RECT 1288.29 599.405 1291.1 618.3 ;
      RECT 1282.67 0 1285.48 37.065 ;
      RECT 1282.67 599.405 1285.48 618.3 ;
      RECT 1243.33 0 1246.14 30.425 ;
      RECT 1243.33 599.405 1246.14 618.3 ;
      RECT 1237.71 0 1240.52 37.065 ;
      RECT 1237.71 599.405 1240.52 618.3 ;
      RECT 1198.37 0 1201.18 30.425 ;
      RECT 1198.37 599.405 1201.18 618.3 ;
      RECT 1192.75 0 1195.56 37.065 ;
      RECT 1192.75 599.405 1195.56 618.3 ;
      RECT 1153.41 0 1156.22 30.425 ;
      RECT 1153.41 599.405 1156.22 618.3 ;
      RECT 1147.79 0 1150.6 37.065 ;
      RECT 1147.79 599.405 1150.6 618.3 ;
      RECT 1108.45 0 1111.26 30.425 ;
      RECT 1108.45 599.405 1111.26 618.3 ;
      RECT 1102.83 0 1105.64 37.065 ;
      RECT 1102.83 599.405 1105.64 618.3 ;
      RECT 1063.49 0 1066.3 30.425 ;
      RECT 1063.49 599.405 1066.3 618.3 ;
      RECT 1057.87 0 1060.68 37.065 ;
      RECT 1057.87 599.405 1060.68 618.3 ;
      RECT 1018.53 0 1021.34 30.425 ;
      RECT 1018.53 599.405 1021.34 618.3 ;
      RECT 1012.91 0 1015.72 37.065 ;
      RECT 1012.91 599.405 1015.72 618.3 ;
      RECT 973.57 0 976.38 30.425 ;
      RECT 973.57 599.405 976.38 618.3 ;
      RECT 967.95 0 970.76 37.065 ;
      RECT 967.95 599.405 970.76 618.3 ;
      RECT 928.61 0 931.42 30.425 ;
      RECT 928.61 599.405 931.42 618.3 ;
      RECT 922.99 0 925.8 37.065 ;
      RECT 922.99 599.405 925.8 618.3 ;
      RECT 883.65 0 886.46 30.425 ;
      RECT 883.65 599.405 886.46 618.3 ;
      RECT 878.03 0 880.84 37.065 ;
      RECT 878.03 599.405 880.84 618.3 ;
      RECT 838.69 0 841.5 30.425 ;
  END
END RM_IHPSG13_1P_8192x32_c4_bm_bist

END LIBRARY
